*** Title:

.include 'translr.net'
.include 'translr.sim'

.model nmos_tkt2.1 nmos level=49 wmax=4e-007 wmin=3e-007 lmax=3e-007 lmin=2.4e-007 version=3.2 mobmod=1 capmod=1 nqsmod=0 binunit=2 binflag=1 tox=5.05e-009 toxm=5.05e-009 xj=1e-007 nch=2.37707e+017 vth0=0.854226 lvth0=-6.45009e-008 
+ wvth0=-2.10231e-007 pvth0=4.41876e-014 vfb=-0.62832 k1=-2.02805 lk1=7.38043e-007 wk1=7.52089e-007 pk1=-2.32679e-013 k2=0.614775 lk2=-1.94265e-007 wk2=-1.91157e-007 pk2=5.69478e-014 k3=0 k3b=0 w0=0 nlx=0 dvt0w=0 dvt1w=0 dvt2w=0 dvt0=0 dvt1=0 dvt2=0 
+ u0=-0.00211838 lu0=8.89274e-009 wu0=1.05834e-008 pu0=-3.24809e-015 ua=-1.80963e-009 lua=-1.36076e-016 wua=9.86002e-016 pua=-5.69659e-023 ub=-5.60906e-018 lub=2.44086e-024 wub=2.04376e-024 pub=-6.21377e-031 uc=-7.98777e-010 luc=2.63925e-016 
+ wuc=2.99104e-016 puc=-8.61043e-023 vsat=62081.5 lvsat=0.00544917 wvsat=0.00575808 pvsat=-2.47655e-009 a0=-3.63456 la0=9.7967e-007 wa0=1.25452e-006 pa0=-3.20869e-013 ags=1.23353 lags=-3.29648e-007 wags=-4.2406e-007 pags=1.13294e-013 b0=0 b1=0 
+ keta=-0.0484089 lketa=1.29448e-008 wketa=1.81329e-008 pketa=-4.24662e-015 a1=0 a2=0.99 rdsw=10 prwg=0.2 prwb=-0.3 wr=1 wint=0 lint=0 dwg=0 dwb=0 voff=-0.631153 lvoff=1.35751e-007 wvoff=1.82641e-007 pvoff=-4.64147e-014 nfactor=-7.09715 
+ lnfactor=1.30782e-006 wnfactor=3.32689e-006 pnfactor=-5.7852e-013 eta0=-0.0169668 leta0=6.83101e-009 weta0=7.24918e-010 peta0=-3.43362e-016 etab=0.0087091 letab=-3.26794e-009 wetab=-3.20679e-009 petab=9.99283e-016 pclm=4.2861 lpclm=-8.1164e-007 
+ wpclm=-1.235e-006 ppclm=2.9187e-013 pdiblc1=0 pdiblc2=0.0892914 lpdiblc2=-2.03446e-008 wpdiblc2=-2.32308e-008 ppdiblc2=6.64669e-015 pdiblcb=-0.0847912 lpdiblcb=1.25288e-007 wpdiblcb=1.21978e-007 ppdiblcb=-5.25336e-014 drout=0 pscbe1=7.70752e+008 
+ pscbe2=1e-020 pvag=0.343793 lpvag=-1.03138e-007 wpvag=-1.37517e-007 ppvag=4.12552e-014 delta=0.01 ngate=1e+030 dsub=0 cit=0.0188351 lcit=-4.10067e-009 wcit=-6.79356e-009 pcit=1.51532e-015 cdsc=0 cdscd=6.21983e-005 lcdscd=-1.95483e-011 
+ wcdscd=-2.48793e-011 pcdscd=7.81931e-018 cdscb=0 xpart=0 cgso=3.15e-010 cgdo=3.15e-010 cgbo=1e-013 cgsl=0 cgdl=0 ckappa=0.6 cf=0 clc=1e-007 cle=0.6 dlc=0 dwc=0 vfbcv=-0.720472 noff=1 voffcv=0 acde=0.5 moin=15 wln=1 wl=0 wwn=1 ww=0 wwl=0 lln=1 ll=0 
+ lwn=1 lw=0 lwl=0 llc=0 lwc=0 lwlc=0 wlc=0 wwc=0 wwlc=0 alpha0=0 alpha1=0 beta0=30 af=1.09369 kf=4.13676e-023 rsh=4 js=0.0001 jsw=0 cj=0.00121101 mj=0.398913 pb=0.786344 cjsw=5.3952e-011 mjsw=2 tref=27 prt=0.628378 ute=-1.29285 kt1=-0.227499 kt1l=0 
+ kt2=-0.0211773 ua1=5.21908e-010 ub1=9.72591e-019 uc1=2.64618e-011 at=10798.4 xti=3 tcj=0.00092022 tcjsw=-0.0079958 tpb=0.0022292 tpbsw=-0.0087143 elm=5 xl=0 xw=0 ldif=1e-007 hdif=2.7e-007 lmlt=1 wmlt=1 rd=0 rdc=0 rs=0 rsc=0 php=0.8 cjgate=2e-014 
+ n=1 

.model nmos_tkt2.2 nmos level=49 wmax=4e-007 wmin=3e-007 lmax=5e-007 lmin=3e-007 acm=2 version=3.2 mobmod=1 capmod=1 nqsmod=0 binunit=2 binflag=1 tox=5.05e-009 toxm=5.05e-009 xj=1e-007 nch=2.37707e+017 vth0=0.658511 lvth0=-5.78649e-009 
+ wvth0=-9.97789e-008 pvth0=1.1052e-014 vfb=-0.62832 k1=1.28389 lk1=-2.5554e-007 wk1=-3.40358e-007 pk1=9.50552e-014 k2=-0.180045 lk2=4.41805e-008 wk2=6.38065e-008 pk2=-1.95411e-014 k3=0 k3b=0 w0=0 nlx=0 dvt0w=0 dvt1w=0 dvt2w=0 dvt0=0 dvt1=0 dvt2=0 
+ u0=0.0452484 lu0=-5.31731e-009 wu0=-1.04058e-008 pu0=3.04869e-015 ua=1.60828e-009 lua=-1.16145e-015 wua=-9.23964e-016 pua=5.16024e-022 ub=1.58318e-018 lub=2.83191e-025 wub=-1.24136e-025 pub=2.89933e-032 uc=2.53e-010 luc=-5.16077e-017 
+ wuc=-1.03666e-016 puc=3.47266e-023 vsat=177278 lvsat=-0.0291098 wvsat=-0.019286 pvsat=5.03668e-009 a0=1.71663 la0=-6.25687e-007 wa0=-2.02329e-007 pa0=1.16185e-013 ags=0.0913679 lags=1.30017e-008 wags=-3.34104e-008 pags=-3.9005e-015 b0=0 b1=0 
+ keta=-0.0526489 lketa=1.42168e-008 wketa=1.53821e-008 pketa=-3.42138e-015 a1=0 a2=0.99 rdsw=10 prwg=0.2 prwb=-0.3 wr=1 wint=0 lint=0 dwg=0 dwb=0 voff=0.0304226 lvoff=-6.27219e-008 wvoff=-6.12641e-008 pvoff=2.67566e-014 nfactor=5.14963 
+ lnfactor=-2.36622e-006 wnfactor=-9.10643e-007 pnfactor=6.92742e-013 eta0=-0.00434049 leta0=3.04311e-009 weta0=-2.25906e-010 peta0=-5.81149e-017 etab=0.00300863 letab=-1.5578e-009 wetab=-1.4973e-010 petab=8.21645e-017 pclm=-1.71178 
+ lpclm=9.87724e-007 wpclm=1.09391e-006 ppclm=-4.06801e-013 pdiblc1=0 pdiblc2=0.0412922 lpdiblc2=-5.94486e-009 wpdiblc2=4.97274e-009 ppdiblc2=-1.81438e-015 pdiblcb=-0.0437246 lpdiblcb=1.12968e-007 wpdiblcb=5.75599e-008 ppdiblcb=-3.32083e-014 drout=0 
+ pscbe1=7.70752e+008 pscbe2=1e-020 pvag=2.5 lpvag=-7.5e-007 delta=0.01 ngate=1e+030 dsub=0 cit=-0.00945375 lcit=4.38599e-009 wcit=2.70651e-009 pcit=-1.3347e-015 cdsc=0 cdscd=-0.000110879 lcdscd=3.23748e-011 wcdscd=4.43514e-011 pcdscd=-1.29499e-017 
+ cdscb=0 xpart=0 cgso=3.15e-010 cgdo=3.15e-010 cgbo=1e-013 cgsl=0 cgdl=0 ckappa=0.6 cf=0 clc=1e-007 cle=0.6 dlc=0 dwc=0 vfbcv=-0.720472 noff=1 voffcv=0 acde=0.5 moin=15 wln=1 wl=0 wwn=1 ww=0 wwl=0 lln=1 ll=0 lwn=1 lw=0 lwl=0 llc=0 lwc=0 lwlc=0 
+ wlc=0 wwc=0 wwlc=0 alpha0=0 alpha1=0 beta0=30 af=1.09369 kf=4.13676e-023 rsh=4 js=0.0001 jsw=0 cj=0.00121101 mj=0.398913 pb=0.786344 cjsw=5.3952e-011 mjsw=2 tref=27 prt=0.628378 ute=-1.29285 kt1=-0.227499 kt1l=0 kt2=-0.0211773 ua1=5.21908e-010 
+ ub1=9.72591e-019 uc1=2.64618e-011 at=10798.4 xti=3 tcj=0.00092022 tcjsw=-0.0079958 tpb=0.0022292 tpbsw=-0.0087143 elm=5 xl=0 xw=0 ldif=1e-007 hdif=2.7e-007 lmlt=1 wmlt=1 rd=0 rdc=0 rs=0 rsc=0 php=0.8 cjgate=2e-014 n=1 

.model nmos_tkt2.3 nmos level=49 wmax=4e-007 wmin=3e-007 lmax=1e-006 lmin=5e-007 acm=2 version=3.2 mobmod=1 capmod=1 nqsmod=0 binunit=2 binflag=1 tox=5.05e-009 toxm=5.05e-009 xj=1e-007 nch=2.37707e+017 vth0=0.481705 lvth0=8.26166e-008 
+ wvth0=-4.62939e-008 pvth0=-1.56905e-014 vfb=-0.62832 k1=0.469168 lk1=1.5182e-007 wk1=-3.60676e-008 pk1=-5.70901e-014 k2=-0.0066459 lk2=-4.25189e-008 wk2=-2.65152e-009 pk2=1.36879e-014 k3=0 k3b=0 w0=0 nlx=0 dvt0w=0 dvt1w=0 dvt2w=0 dvt0=0 dvt1=0 
+ dvt2=0 u0=0.0344002 lu0=1.06798e-010 wu0=-3.80659e-009 pu0=-2.5093e-016 ua=-1.18702e-010 lua=-2.97957e-016 wua=1.25576e-018 pua=5.34139e-023 ub=1.14852e-018 lub=5.00524e-025 wub=5.70785e-026 pub=-6.16137e-032 uc=6.48153e-011 luc=4.24845e-017 
+ wuc=-2.45795e-017 puc=-4.81666e-024 vsat=880942 lvsat=-0.380942 wvsat=0.00921266 pvsat=-9.21267e-009 a0=2.5023 la0=-1.01852e-006 wa0=-2.27904e-007 pa0=1.28973e-013 ags=-0.0773712 lags=9.73712e-008 wags=4.12114e-008 pags=-4.12114e-014 b0=0 b1=0 
+ keta=0.0872715 lketa=-5.57434e-008 wketa=-2.18284e-008 pketa=1.51839e-014 a1=0 a2=0.99 rdsw=10 prwg=0.2 prwb=-0.3 wr=1 wint=0 lint=0 dwg=0 dwb=0 voff=-0.106527 lvoff=5.75279e-009 wvoff=5.75591e-009 pvoff=-6.75336e-015 nfactor=-7.12917 
+ lnfactor=3.77319e-006 wnfactor=2.73875e-006 pnfactor=-1.13196e-012 eta0=0.0132777 leta0=-5.766e-009 weta0=-3.68401e-009 peta0=1.67094e-015 etab=0.000106965 letab=-1.06965e-010 wetab=-1.45986e-011 petab=1.45986e-017 pclm=-13.9359 lpclm=7.0998e-006 
+ wpclm=6.82138e-006 ppclm=-3.27054e-012 pdiblc1=0 pdiblc2=-0.529978 lpdiblc2=2.7969e-007 wpdiblc2=2.08829e-007 ppdiblc2=-1.03742e-013 pdiblcb=2.61779 lpdiblcb=-1.21779e-006 wpdiblcb=-9.51143e-007 ppdiblcb=4.71143e-013 drout=0 pscbe1=7.70752e+008 
+ pscbe2=1e-020 pvag=7 lpvag=-3e-006 wpvag=-2.4e-006 ppvag=1.2e-012 delta=0.01 ngate=1e+030 dsub=0 cit=0.00753132 lcit=-4.10654e-009 wcit=-2.58429e-009 pcit=1.3107e-015 cdsc=0 cdscd=1.15393e-005 lcdscd=-2.88342e-011 wcdscd=-4.61573e-012 
+ pcdscd=1.15337e-017 cdscb=0 xpart=0 cgso=3.15e-010 cgdo=3.15e-010 cgbo=1e-013 cgsl=0 cgdl=0 ckappa=0.6 cf=0 clc=1e-007 cle=0.6 dlc=0 dwc=0 vfbcv=-0.720472 noff=1 voffcv=0 acde=0.5 moin=15 wln=1 wl=0 wwn=1 ww=0 wwl=0 lln=1 ll=0 lwn=1 lw=0 lwl=0 
+ llc=0 lwc=0 lwlc=0 wlc=0 wwc=0 wwlc=0 alpha0=0 alpha1=0 beta0=30 af=1.09369 kf=4.13676e-023 rsh=4 js=0.0001 jsw=0 cj=0.00121101 mj=0.398913 pb=0.786344 cjsw=5.3952e-011 mjsw=2 tref=27 prt=0.628378 ute=-1.29285 kt1=-0.227499 kt1l=0 kt2=-0.0211773 
+ ua1=5.21908e-010 ub1=9.72591e-019 uc1=2.64618e-011 at=10798.4 xti=3 tcj=0.00092022 tcjsw=-0.0079958 tpb=0.0022292 tpbsw=-0.0087143 elm=5 xl=0 xw=0 ldif=1e-007 hdif=2.7e-007 lmlt=1 wmlt=1 rd=0 rdc=0 rs=0 rsc=0 php=0.8 cjgate=2e-014 n=1 

.model nmos_tkt2.4 nmos level=49 wmax=4e-007 wmin=3e-007 lmax=1e-005 lmin=1e-006 acm=2 version=3.2 mobmod=1 capmod=1 nqsmod=0 binunit=2 binflag=1 tox=5.05e-009 toxm=5.05e-009 xj=1e-007 nch=2.37707e+017 vth0=0.482813 lvth0=8.1509e-008 
+ wvth0=-5.94361e-008 pvth0=-2.54826e-015 vfb=-0.62832 k1=0.447189 lk1=1.73799e-007 wk1=-1.99638e-008 pk1=-7.31939e-014 k2=0.0218474 lk2=-7.10122e-008 wk2=-1.30074e-008 pk2=2.40438e-014 k3=0 k3b=0 w0=0 nlx=0 dvt0w=0 dvt1w=0 dvt2w=0 dvt0=0 dvt1=0 
+ dvt2=0 u0=0.0327944 lu0=1.71258e-009 wu0=-3.78262e-009 pu0=-2.749e-016 ua=-5.64417e-010 lua=1.47758e-016 wua=1.32915e-016 pua=-7.82451e-023 ub=1.51716e-018 lub=1.31884e-025 wub=-8.24053e-026 pub=7.78701e-032 uc=4.30165e-011 luc=6.42833e-017 
+ wuc=-2.04235e-017 puc=-8.9727e-024 vsat=500000 a0=0.756867 la0=7.26908e-007 wa0=-1.25702e-007 pa0=2.67708e-014 ags=0.02 b0=0 b1=0 keta=0.0120957 lketa=1.94324e-008 wketa=-7.89781e-010 pketa=-5.85476e-015 a1=0 a2=0.99 rdsw=10 prwg=0.2 prwb=-0.3 
+ wr=1 wint=0 lint=0 dwg=0 dwb=0 voff=-0.166132 lvoff=6.53577e-008 wvoff=2.06721e-008 pvoff=-2.16695e-014 nfactor=-0.686862 lnfactor=-2.66912e-006 wnfactor=2.45367e-007 pnfactor=1.36143e-012 eta0=0.00112498 leta0=6.38674e-009 weta0=-2.32878e-010 
+ peta0=-1.7802e-015 etab=0 pclm=6.31513 lpclm=-1.31513e-005 wpclm=-3.94537e-007 ppclm=3.94538e-012 pdiblc1=0 pdiblc2=0.138921 lpdiblc2=-3.89209e-007 wpdiblc2=-1.16763e-008 ppdiblc2=1.16763e-013 pdiblcb=0.0666665 lpdiblcb=1.33333e-006 
+ wpdiblcb=5.33333e-008 ppdiblcb=-5.33333e-013 drout=0 pscbe1=7.70752e+008 pscbe2=1e-020 pvag=-0.444445 lpvag=4.44444e-006 wpvag=1.33333e-007 ppvag=-1.33333e-012 delta=0.01 ngate=1e+030 dsub=0 cit=-2.09521e-005 lcit=3.44572e-009 wcit=1.94209e-011 
+ pcit=-1.29301e-015 cdsc=0 cdscd=7.52641e-005 lcdscd=-9.2559e-011 wcdscd=-2.27714e-011 pcdscd=2.96893e-017 cdscb=0 xpart=0 cgso=3.15e-010 cgdo=3.15e-010 cgbo=1e-013 cgsl=0 cgdl=0 ckappa=0.6 cf=0 clc=1e-007 cle=0.6 dlc=0 dwc=0 vfbcv=-0.720472 noff=1 
+ voffcv=0 acde=0.5 moin=15 wln=1 wl=0 wwn=1 ww=0 wwl=0 lln=1 ll=0 lwn=1 lw=0 lwl=0 llc=0 lwc=0 lwlc=0 wlc=0 wwc=0 wwlc=0 alpha0=0 alpha1=0 beta0=30 af=1.09369 kf=4.13676e-023 rsh=4 js=0.0001 jsw=0 cj=0.00121101 mj=0.398913 pb=0.786344 
+ cjsw=5.3952e-011 mjsw=2 tref=27 prt=0.628378 ute=-1.29285 kt1=-0.227499 kt1l=0 kt2=-0.0211773 ua1=5.21908e-010 ub1=9.72591e-019 uc1=2.64618e-011 at=10798.4 xti=3 tcj=0.00092022 tcjsw=-0.0079958 tpb=0.0022292 tpbsw=-0.0087143 elm=5 xl=0 xw=0 
+ ldif=1e-007 hdif=2.7e-007 lmlt=1 wmlt=1 rd=0 rdc=0 rs=0 rsc=0 php=0.8 cjgate=2e-014 n=1 

.model nmos_tkt2.5 nmos level=49 wmax=4e-007 wmin=3e-007 lmax=2e-005 lmin=1e-005 acm=2 version=3.2 mobmod=1 capmod=1 nqsmod=0 binunit=2 binflag=1 tox=5.05e-009 toxm=5.05e-009 xj=1e-007 nch=2.37707e+017 vth0=0.490964 wvth0=-5.96909e-008 vfb=-0.62832 
+ k1=0.464569 wk1=-2.72832e-008 k2=0.0147462 wk2=-1.0603e-008 k3=0 k3b=0 w0=0 nlx=0 dvt0w=0 dvt1w=0 dvt2w=0 dvt0=0 dvt1=0 dvt2=0 u0=0.0329657 wu0=-3.8101e-009 ua=-5.49641e-010 wua=1.2509e-016 ub=1.53035e-018 wub=-7.46183e-026 uc=4.94448e-011 
+ wuc=-2.13208e-017 vsat=500000 a0=0.829557 wa0=-1.23025e-007 ags=0.02 b0=0 b1=0 keta=0.014039 wketa=-1.37526e-009 a1=0 a2=0.99 rdsw=10 prwg=0.2 prwb=-0.3 wr=1 wint=0 lint=0 dwg=0 dwb=0 voff=-0.159596 wvoff=1.85051e-008 nfactor=-0.953775 
+ wnfactor=3.8151e-007 eta0=0.00176365 weta0=-4.10897e-010 etab=0 pclm=5 pdiblc1=0 pdiblc2=0.1 pdiblcb=0.2 drout=0 pscbe1=7.70752e+008 pscbe2=1e-020 pvag=0 delta=0.01 ngate=1e+030 dsub=0 cit=0.000323621 wcit=-1.0988e-010 cdsc=0 cdscd=6.60082e-005 
+ wcdscd=-1.98025e-011 cdscb=0 xpart=0 cgso=3.15e-010 cgdo=3.15e-010 cgbo=1e-013 cgsl=0 cgdl=0 ckappa=0.6 cf=0 clc=1e-007 cle=0.6 dlc=0 dwc=0 vfbcv=-0.720472 noff=1 voffcv=0 acde=0.5 moin=15 wln=1 wl=0 wwn=1 ww=0 wwl=0 lln=1 ll=0 lwn=1 lw=0 lwl=0 
+ llc=0 lwc=0 lwlc=0 wlc=0 wwc=0 wwlc=0 alpha0=0 alpha1=0 beta0=30 af=1.09369 kf=4.13676e-023 rsh=4 js=0.0001 jsw=0 cj=0.00121101 mj=0.398913 pb=0.786344 cjsw=5.3952e-011 mjsw=2 tref=27 prt=0.628378 ute=-1.29285 kt1=-0.227499 kt1l=0 kt2=-0.0211773 
+ ua1=5.21908e-010 ub1=9.72591e-019 uc1=2.64618e-011 at=10798.4 xti=3 tcj=0.00092022 tcjsw=-0.0079958 tpb=0.0022292 tpbsw=-0.0087143 elm=5 xl=0 xw=0 ldif=1e-007 hdif=2.7e-007 lmlt=1 wmlt=1 rd=0 rdc=0 rs=0 rsc=0 php=0.8 cjgate=2e-014 n=1 

.model nmos_tkt2.6 nmos level=49 wmax=1e-006 wmin=4e-007 lmax=3e-007 lmin=2.4e-007 acm=2 version=3.2 mobmod=1 capmod=1 nqsmod=0 binunit=2 binflag=1 tox=5.05e-009 toxm=5.05e-009 xj=1e-007 nch=2.37707e+017 vth0=0.32427 lvth0=6.90065e-008 
+ wvth0=1.75173e-009 pvth0=-9.2154e-015 vfb=-0.62832 k1=1.09162 lk1=-1.09725e-007 wk1=-4.95781e-007 pk1=1.06428e-013 k2=-0.157401 lk2=1.08138e-008 wk2=1.17714e-007 pk2=-2.50839e-014 k3=0 k3b=0 w0=0 nlx=0 dvt0w=0 dvt1w=0 dvt2w=0 dvt0=0 dvt1=0 dvt2=0 
+ u0=0.0359344 lu0=1.95269e-010 wu0=-4.63766e-009 pu0=2.30898e-016 ua=-1.27858e-009 lua=1.8566e-016 wua=7.73584e-016 pua=-1.8566e-022 ub=3.45618e-018 lub=-1.40065e-025 wub=-1.58233e-024 pub=4.10995e-031 uc=3.0603e-010 luc=-3.1166e-017 
+ wuc=-1.42819e-016 puc=3.19322e-023 vsat=79350.4 lvsat=-0.000565897 wvsat=-0.00114949 pvsat=-7.0525e-011 a0=0.607702 la0=-2.24457e-007 wa0=-4.42386e-007 pa0=1.60782e-013 ags=-0.111794 lags=3.80305e-008 wags=1.14071e-007 pags=-3.3777e-014 b0=0 b1=0 
+ keta=0.0158994 lketa=-9.44393e-009 wketa=-7.59041e-009 pketa=4.70886e-015 a1=0 a2=0.99 rdsw=10 prwg=0.2 prwb=-0.3 wr=1 wint=0 lint=0 dwg=0 dwb=0 voff=0.214534 lvoff=-9.2244e-008 wvoff=-1.55634e-007 pvoff=4.47832e-014 nfactor=-2.46119 
+ lnfactor=6.31503e-007 wnfactor=1.47251e-006 pnfactor=-3.07994e-013 eta0=0.00388266 leta0=4.14113e-010 weta0=-7.61488e-009 peta0=2.2234e-015 etab=0.00109705 letab=-9.73671e-010 wetab=-1.61973e-010 petab=8.1576e-017 pclm=-0.38818 lpclm=4.36774e-007 
+ wpclm=6.34716e-007 ppclm=-2.07496e-013 pdiblc1=0 pdiblc2=-0.0749098 lpdiblc2=2.6653e-008 wpdiblc2=4.24497e-008 ppdiblc2=-1.21523e-014 pdiblcb=0.391929 lpdiblcb=-1.33605e-007 wpdiblcb=-6.87101e-008 ppdiblcb=5.10236e-014 drout=0 pscbe1=7.70752e+008 
+ pscbe2=1e-020 pvag=-0.666239 lpvag=1.99872e-007 wpvag=2.66496e-007 ppvag=-7.99488e-014 delta=0.01 ngate=1e+030 dsub=0 cit=0.00446295 lcit=-8.27478e-010 wcit=-1.0447e-009 pcit=2.06043e-016 cdsc=0 cdscd=-9.09851e-005 lcdscd=2.72955e-011 
+ wcdscd=3.6394e-011 pcdscd=-1.09182e-017 cdscb=0 xpart=0 cgso=3.15e-010 cgdo=3.15e-010 cgbo=1e-013 cgsl=0 cgdl=0 ckappa=0.6 cf=0 clc=1e-007 cle=0.6 dlc=0 dwc=0 vfbcv=-0.720472 noff=1 voffcv=0 acde=0.5 moin=15 wln=1 wl=0 wwn=1 ww=0 wwl=0 lln=1 ll=0 
+ lwn=1 lw=0 lwl=0 llc=0 lwc=0 lwlc=0 wlc=0 wwc=0 wwlc=0 alpha0=0 alpha1=0 beta0=30 af=1.09369 kf=4.13676e-023 rsh=4 js=0.0001 jsw=0 cj=0.00121101 mj=0.398913 pb=0.786344 cjsw=5.3952e-011 mjsw=2 tref=27 prt=0.628378 ute=-1.29285 kt1=-0.227499 kt1l=0 
+ kt2=-0.0211773 ua1=5.21908e-010 ub1=9.72591e-019 uc1=2.64618e-011 at=10798.4 xti=3 tcj=0.00092022 tcjsw=-0.0079958 tpb=0.0022292 tpbsw=-0.0087143 elm=5 xl=0 xw=0 ldif=1e-007 hdif=2.7e-007 lmlt=1 wmlt=1 rd=0 rdc=0 rs=0 rsc=0 php=0.8 cjgate=2e-014 
+ n=1 

.model nmos_tkt2.7 nmos level=49 wmax=1e-006 wmin=4e-007 lmax=5e-007 lmin=3e-007 acm=2 version=3.2 mobmod=1 capmod=1 nqsmod=0 binunit=2 binflag=1 tox=5.05e-009 toxm=5.05e-009 xj=1e-007 nch=2.37707e+017 vth0=0.482646 lvth0=2.14937e-008 
+ wvth0=-2.94328e-008 pvth0=1.39952e-016 vfb=-0.62832 k1=0.197629 lk1=1.58473e-007 wk1=9.4145e-008 pk1=-7.05499e-014 k2=0.104084 lk2=-6.76317e-008 wk2=-4.9845e-008 pk2=2.51838e-014 k3=0 k3b=0 w0=0 nlx=0 dvt0w=0 dvt1w=0 dvt2w=0 dvt0=0 dvt1=0 dvt2=0 
+ u0=0.0327943 lu0=1.13729e-009 wu0=-5.42418e-009 pu0=4.66854e-016 ua=-3.73913e-010 lua=-8.57412e-017 wua=-1.31087e-016 pua=8.57412e-023 ub=1.33699e-018 lub=4.95692e-025 wub=-2.56585e-026 pub=-5.60069e-032 uc=6.71612e-011 luc=4.04948e-017 
+ wuc=-2.93306e-017 puc=-2.1144e-024 vsat=123826 lvsat=-0.0139086 wvsat=0.00209474 pvsat=-1.0438e-009 a0=1.80278 la0=-5.82981e-007 wa0=-2.36791e-007 pa0=9.91029e-014 ags=-0.0153352 lags=9.09292e-009 wags=9.27086e-009 pags=-2.337e-015 b0=0 b1=0 
+ keta=0.0232393 lketa=-1.16459e-008 wketa=-1.49732e-008 pketa=6.92369e-015 a1=0 a2=0.99 rdsw=10 prwg=0.2 prwb=-0.3 wr=1 wint=0 lint=0 dwg=0 dwb=0 voff=-0.207465 lvoff=3.43556e-008 wvoff=3.38909e-008 pvoff=-1.20744e-014 nfactor=-2.13955 
+ lnfactor=5.35011e-007 wnfactor=2.00503e-006 pnfactor=-4.67749e-013 eta0=1.42008e-005 leta0=1.57465e-009 weta0=-1.96778e-009 peta0=5.29267e-016 etab=0.000400752 letab=-7.64781e-010 wetab=8.93422e-010 petab=-2.35042e-016 pclm=0.6598 
+ lpclm=1.2238e-007 wpclm=1.45274e-007 ppclm=-6.06629e-014 pdiblc1=0 pdiblc2=-0.0136541 lpdiblc2=8.27624e-009 wpdiblc2=2.69513e-008 ppdiblc2=-7.50281e-015 pdiblcb=0.0827491 lpdiblcb=-4.08512e-008 wpdiblcb=6.97036e-009 ppdiblcb=2.83195e-014 drout=0 
+ pscbe1=7.70752e+008 pscbe2=1e-020 pvag=1.06228 lpvag=-3.18683e-007 wpvag=5.7509e-007 ppvag=-1.72527e-013 delta=0.01 ngate=1e+030 dsub=0 cit=0.00455528 lcit=-8.55175e-010 wcit=-2.8971e-009 pcit=7.61762e-016 cdsc=0 cdscd=0 cdscb=0 xpart=0 
+ cgso=3.15e-010 cgdo=3.15e-010 cgbo=1e-013 cgsl=0 cgdl=0 ckappa=0.6 cf=0 clc=1e-007 cle=0.6 dlc=0 dwc=0 vfbcv=-0.720472 noff=1 voffcv=0 acde=0.5 moin=15 wln=1 wl=0 wwn=1 ww=0 wwl=0 lln=1 ll=0 lwn=1 lw=0 lwl=0 llc=0 lwc=0 lwlc=0 wlc=0 wwc=0 wwlc=0 
+ alpha0=0 alpha1=0 beta0=30 af=1.09369 kf=4.13676e-023 rsh=4 js=0.0001 jsw=0 cj=0.00121101 mj=0.398913 pb=0.786344 cjsw=5.3952e-011 mjsw=2 tref=27 prt=0.628378 ute=-1.29285 kt1=-0.227499 kt1l=0 kt2=-0.0211773 ua1=5.21908e-010 ub1=9.72591e-019 
+ uc1=2.64618e-011 at=10798.4 xti=3 tcj=0.00092022 tcjsw=-0.0079958 tpb=0.0022292 tpbsw=-0.0087143 elm=5 xl=0 xw=0 ldif=1e-007 hdif=2.7e-007 lmlt=1 wmlt=1 rd=0 rdc=0 rs=0 rsc=0 php=0.8 cjgate=2e-014 n=1 

.model nmos_tkt2.8 nmos level=49 wmax=1e-006 wmin=4e-007 lmax=1e-006 lmin=5e-007 acm=2 version=3.2 mobmod=1 capmod=1 nqsmod=0 binunit=2 binflag=1 tox=5.05e-009 toxm=5.05e-009 xj=1e-007 nch=2.37707e+017 vth0=0.446967 lvth0=3.93335e-008 
+ wvth0=-3.23985e-008 pvth0=1.6228e-015 vfb=-0.62832 k1=0.343737 lk1=8.54195e-008 wk1=1.41051e-008 pk1=-3.053e-014 k2=0.0348105 lk2=-3.2995e-008 wk2=-1.92341e-008 pk2=9.87834e-015 k3=0 k3b=0 w0=0 nlx=0 dvt0w=0 dvt1w=0 dvt2w=0 dvt0=0 dvt1=0 dvt2=0 
+ u0=0.0277163 lu0=3.67627e-009 wu0=-1.13303e-009 pu0=-1.67872e-015 ua=-7.64625e-010 lua=1.09615e-016 wua=2.59625e-016 pua=-1.09615e-022 ub=1.54347e-018 lub=3.92451e-025 wub=-1.00903e-025 pub=-1.83848e-032 uc=8.25081e-012 luc=6.995e-017 
+ wuc=-1.95374e-018 puc=-1.58028e-023 vsat=903991 lvsat=-0.403991 pvsat=7.15104e-012 a0=1.55942 la0=-4.61301e-007 wa0=1.49247e-007 pa0=-9.39156e-014 ags=-0.096184 lags=4.95173e-008 wags=4.87365e-008 pags=-2.20698e-014 b0=0 b1=0 keta=0.0103598 
+ lketa=-5.20614e-009 wketa=8.93625e-009 pketa=-5.03102e-015 a1=0 a2=0.99 rdsw=10 prwg=0.2 prwb=-0.3 wr=1 wint=0 lint=0 dwg=0 dwb=0 voff=-0.160783 lvoff=1.10146e-008 wvoff=2.74583e-008 pvoff=-8.85806e-015 nfactor=0.188195 lnfactor=-6.28864e-007 
+ wnfactor=-1.88195e-007 pnfactor=6.28864e-013 eta0=-0.00499448 leta0=4.07899e-009 weta0=3.62487e-009 peta0=-2.26706e-015 etab=0.000721124 letab=-9.24967e-010 wetab=-2.60262e-010 petab=3.41799e-016 pclm=13.0408 lpclm=-6.06813e-006 
+ wpclm=-3.96933e-006 ppclm=1.99664e-012 pdiblc1=0 pdiblc2=0.313864 lpdiblc2=-1.55483e-007 wpdiblc2=-1.28708e-007 ppdiblc2=7.03269e-014 pdiblcb=0.398953 lpdiblcb=-1.98953e-007 wpdiblcb=-6.36093e-008 ppdiblcb=6.36093e-014 drout=0 pscbe1=7.70752e+008 
+ pscbe2=1e-020 pvag=-1.75824 lpvag=1.09158e-006 wpvag=1.1033e-006 ppvag=-4.36631e-013 delta=0.01 ngate=1e+030 dsub=0 cit=-0.000532847 lcit=1.68889e-009 wcit=6.41373e-010 pcit=-1.00747e-015 cdsc=0 cdscd=0.000126572 lcdscd=-6.32861e-011 
+ wcdscd=-5.06289e-011 pcdscd=2.53145e-017 cdscb=0 xpart=0 cgso=3.15e-010 cgdo=3.15e-010 cgbo=1e-013 cgsl=0 cgdl=0 ckappa=0.6 cf=0 clc=1e-007 cle=0.6 dlc=0 dwc=0 vfbcv=-0.720472 noff=1 voffcv=0 acde=0.5 moin=15 wln=1 wl=0 wwn=1 ww=0 wwl=0 lln=1 ll=0 
+ lwn=1 lw=0 lwl=0 llc=0 lwc=0 lwlc=0 wlc=0 wwc=0 wwlc=0 alpha0=0 alpha1=0 beta0=30 af=1.09369 kf=4.13676e-023 rsh=4 js=0.0001 jsw=0 cj=0.00121101 mj=0.398913 pb=0.786344 cjsw=5.3952e-011 mjsw=2 tref=27 prt=0.628378 ute=-1.29285 kt1=-0.227499 kt1l=0 
+ kt2=-0.0211773 ua1=5.21908e-010 ub1=9.72591e-019 uc1=2.64618e-011 at=10798.4 xti=3 tcj=0.00092022 tcjsw=-0.0079958 tpb=0.0022292 tpbsw=-0.0087143 elm=5 xl=0 xw=0 ldif=1e-007 hdif=2.7e-007 lmlt=1 wmlt=1 rd=0 rdc=0 rs=0 rsc=0 php=0.8 cjgate=2e-014 
+ n=1 

.model nmos_tkt2.9 nmos level=49 wmax=1e-006 wmin=4e-007 lmax=1e-005 lmin=1e-006 acm=2 version=3.2 mobmod=1 capmod=1 nqsmod=0 binunit=2 binflag=1 tox=5.05e-009 toxm=5.05e-009 xj=1e-007 nch=2.37707e+017 vth0=0.419634 lvth0=6.66658e-008 
+ wvth0=-3.41647e-008 pvth0=3.38903e-015 vfb=-0.62832 k1=0.43538 lk1=-6.22404e-009 wk1=-1.52403e-008 pk1=-1.18452e-015 k2=0.00643675 lk2=-4.62125e-009 wk2=-6.84313e-009 pk2=-2.51259e-015 k3=0 k3b=0 w0=0 nlx=0 dvt0w=0 dvt1w=0 dvt2w=0 dvt0=0 dvt1=0 
+ dvt2=0 u0=0.0296864 lu0=1.70622e-009 wu0=-2.53939e-009 pu0=-2.72356e-016 ua=-6.86868e-010 lua=3.18578e-017 wua=1.81895e-016 pua=-3.1885e-023 ub=1.7007e-018 lub=2.35223e-025 wub=-1.55822e-025 pub=3.65347e-032 uc=3.57503e-011 luc=4.24505e-017 
+ wuc=-1.7517e-017 puc=-2.39563e-025 vsat=500000 a0=0.559608 la0=5.38512e-007 wa0=-4.67985e-008 pa0=1.02129e-013 ags=0.0274074 lags=-7.40741e-008 wags=-2.96296e-009 pags=2.96296e-014 b0=0 b1=0 keta=0.0111648 lketa=-6.01112e-009 wketa=-4.17412e-010 
+ pketa=4.32264e-015 a1=0 a2=0.99 rdsw=10 prwg=0.2 prwb=-0.3 wr=1 wint=0 lint=0 dwg=0 dwb=0 voff=-0.149749 lvoff=-1.87025e-011 wvoff=1.41192e-008 pvoff=4.48104e-015 nfactor=0.0489631 lnfactor=-4.89632e-007 wnfactor=-4.89632e-008 
+ pnfactor=4.89632e-013 eta0=0.000208109 leta0=-1.1236e-009 weta0=1.3387e-010 peta0=1.22394e-015 etab=2.26493e-005 letab=-2.26493e-010 wetab=-9.05969e-012 petab=9.0597e-017 pclm=4.78081 lpclm=2.19188e-006 wpclm=2.19188e-007 ppclm=-2.19188e-012 
+ pdiblc1=0 pdiblc2=0.0935132 lpdiblc2=6.48681e-008 wpdiblc2=6.4868e-009 ppdiblc2=-6.48681e-014 pdiblcb=0.2 drout=0 pscbe1=7.70752e+008 pscbe2=1e-020 pvag=0.074074 lpvag=-7.40741e-007 wpvag=-7.4074e-008 ppvag=7.40741e-013 delta=0.01 ngate=1e+030 
+ dsub=0 cit=0.00164245 lcit=-4.86407e-010 wcit=-6.45939e-010 pcit=2.79838e-016 cdsc=0 cdscd=-1.92555e-005 lcdscd=8.25417e-011 wcdscd=1.50365e-011 pcdscd=-4.03509e-017 cdscb=0 xpart=0 cgso=3.15e-010 cgdo=3.15e-010 cgbo=1e-013 cgsl=0 cgdl=0 
+ ckappa=0.6 cf=0 clc=1e-007 cle=0.6 dlc=0 dwc=0 vfbcv=-0.720472 noff=1 voffcv=0 acde=0.5 moin=15 wln=1 wl=0 wwn=1 ww=0 wwl=0 lln=1 ll=0 lwn=1 lw=0 lwl=0 llc=0 lwc=0 lwlc=0 wlc=0 wwc=0 wwlc=0 alpha0=0 alpha1=0 beta0=30 af=1.09369 kf=4.13676e-023 
+ rsh=4 js=0.0001 jsw=0 cj=0.00121101 mj=0.398913 pb=0.786344 cjsw=5.3952e-011 mjsw=2 tref=27 prt=0.628378 ute=-1.29285 kt1=-0.227499 kt1l=0 kt2=-0.0211773 ua1=5.21908e-010 ub1=9.72591e-019 uc1=2.64618e-011 at=10798.4 xti=3 tcj=0.00092022 
+ tcjsw=-0.0079958 tpb=0.0022292 tpbsw=-0.0087143 elm=5 xl=0 xw=0 ldif=1e-007 hdif=2.7e-007 lmlt=1 wmlt=1 rd=0 rdc=0 rs=0 rsc=0 php=0.8 cjgate=2e-014 n=1 

.model nmos_tkt2.10 nmos level=49 wmax=1e-006 wmin=4e-007 lmax=2e-005 lmin=1e-005 acm=2 version=3.2 mobmod=1 capmod=1 nqsmod=0 binunit=2 binflag=1 tox=5.05e-009 toxm=5.05e-009 xj=1e-007 nch=2.37707e+017 vth0=0.426301 wvth0=-3.38258e-008 vfb=-0.62832 
+ k1=0.434758 wk1=-1.53588e-008 k2=0.00597463 wk2=-7.09439e-009 k3=0 k3b=0 w0=0 nlx=0 dvt0w=0 dvt1w=0 dvt2w=0 dvt0=0 dvt1=0 dvt2=0 u0=0.029857 wu0=-2.56663e-009 ua=-6.83682e-010 wua=1.78707e-016 ub=1.72422e-018 wub=-1.52169e-025 uc=3.99954e-011 
+ wuc=-1.7541e-017 vsat=500000 a0=0.613459 wa0=-3.65855e-008 ags=0.02 b0=0 b1=0 keta=0.0105637 wketa=1.48515e-011 a1=0 a2=0.99 rdsw=10 prwg=0.2 prwb=-0.3 wr=1 wint=0 lint=0 dwg=0 dwb=0 voff=-0.149751 wvoff=1.45673e-008 nfactor=0 eta0=9.57488e-005 
+ weta0=2.56264e-010 etab=0 pclm=5 pdiblc1=0 pdiblc2=0.1 pdiblcb=0.2 drout=0 pscbe1=7.70752e+008 pscbe2=1e-020 pvag=0 delta=0.01 ngate=1e+030 dsub=0 cit=0.00159381 wcit=-6.17955e-010 cdsc=0 cdscd=-1.10014e-005 wcdscd=1.10014e-011 cdscb=0 xpart=0 
+ cgso=3.15e-010 cgdo=3.15e-010 cgbo=1e-013 cgsl=0 cgdl=0 ckappa=0.6 cf=0 clc=1e-007 cle=0.6 dlc=0 dwc=0 vfbcv=-0.720472 noff=1 voffcv=0 acde=0.5 moin=15 wln=1 wl=0 wwn=1 ww=0 wwl=0 lln=1 ll=0 lwn=1 lw=0 lwl=0 llc=0 lwc=0 lwlc=0 wlc=0 wwc=0 wwlc=0 
+ alpha0=0 alpha1=0 beta0=30 af=1.09369 kf=4.13676e-023 rsh=4 js=0.0001 jsw=0 cj=0.00121101 mj=0.398913 pb=0.786344 cjsw=5.3952e-011 mjsw=2 tref=27 prt=0.628378 ute=-1.29285 kt1=-0.227499 kt1l=0 kt2=-0.0211773 ua1=5.21908e-010 ub1=9.72591e-019 
+ uc1=2.64618e-011 at=10798.4 xti=3 tcj=0.00092022 tcjsw=-0.0079958 tpb=0.0022292 tpbsw=-0.0087143 elm=5 xl=0 xw=0 ldif=1e-007 hdif=2.7e-007 lmlt=1 wmlt=1 rd=0 rdc=0 rs=0 rsc=0 php=0.8 cjgate=2e-014 n=1 

.model nmos_tkt2.11 nmos level=49 wmax=1e-005 wmin=1e-006 lmax=3e-007 lmin=2.4e-007 acm=2 version=3.2 mobmod=1 capmod=1 nqsmod=0 binunit=2 binflag=1 tox=5.05e-009 toxm=5.05e-009 xj=1e-007 nch=2.37707e+017 vth0=0.546928 lvth0=-1.13902e-009 
+ wvth0=-2.20907e-007 pvth0=6.09302e-014 vfb=-0.62832 k1=0.756508 lk1=-4.73433e-008 wk1=-1.60665e-007 pk1=4.40462e-014 k2=-0.020226 lk2=-1.79222e-008 wk2=-1.9461e-008 pk2=3.65212e-015 k3=0 k3b=0 w0=0 nlx=0 dvt0w=0 dvt1w=0 dvt2w=0 dvt0=0 dvt1=0 
+ dvt2=0 u0=-0.0757849 lu0=3.52419e-008 wu0=1.07082e-007 pu0=-3.48157e-014 ua=-1.0168e-008 lua=2.8989e-015 wua=9.663e-015 pua=-2.8989e-021 ub=-3.00248e-019 lub=1.15184e-024 wub=2.1741e-024 pub=-8.8091e-031 uc=-5.23219e-010 luc=2.28412e-016 
+ wuc=6.8643e-016 puc=-2.27646e-022 vsat=87413.2 lvsat=-0.00177043 wvsat=-0.00921225 pvsat=1.13401e-009 a0=0.657188 la0=-1.68655e-007 wa0=-4.91872e-007 pa0=1.04979e-013 ags=0.0961399 lags=-2.41732e-008 wags=-9.38628e-008 pags=2.84267e-014 b0=0 b1=0 
+ keta=-0.0315879 lketa=7.11274e-009 wketa=3.98969e-008 pketa=-1.18478e-014 a1=0 a2=0.99 rdsw=10 prwg=1.97778 lprwg=-5.33333e-007 wprwg=-1.77778e-006 pprwg=5.33333e-013 prwb=-2.96667 lprwb=8e-007 wprwb=2.66667e-006 pprwb=-8e-013 wr=1 wint=0 lint=0 
+ dwg=0 dwb=0 voff=-0.0660015 lvoff=-7.27479e-009 wvoff=1.24901e-007 pvoff=-4.01861e-014 nfactor=3.11512 lnfactor=-6.70648e-007 wnfactor=-4.1038e-006 pnfactor=9.94157e-013 eta0=-0.0163923 leta0=6.05196e-009 weta0=1.26601e-008 peta0=-3.41445e-015 
+ etab=0.00127062 letab=-1.12312e-009 wetab=-3.35546e-010 petab=2.31028e-016 pclm=0.626383 lpclm=1.93275e-007 wpclm=-3.79847e-007 ppclm=3.60036e-014 pdiblc1=0 pdiblc2=0.0122803 lpdiblc2=3.67442e-009 wpdiblc2=-4.47404e-008 ppdiblc2=1.08262e-014 
+ pdiblcb=-0.381154 lpdiblcb=1.20929e-007 wpdiblcb=7.04373e-007 ppdiblcb=-2.0351e-013 drout=0 pscbe1=7.70752e+008 pscbe2=1e-020 pvag=0.441962 lpvag=4.36119e-008 wpvag=-8.41705e-007 ppvag=7.63112e-014 delta=0.01 ngate=1e+030 dsub=0 cit=-0.00359522 
+ lcit=1.16201e-009 wcit=7.01347e-009 pcit=-1.78344e-015 cdsc=0 cdscd=-0.000177097 lcdscd=5.31291e-011 wcdscd=1.22506e-010 pcdscd=-3.67518e-017 cdscb=0 xpart=0 cgso=3.15e-010 cgdo=3.15e-010 cgbo=1e-013 cgsl=0 cgdl=0 ckappa=0.6 cf=0 clc=1e-007 
+ cle=0.6 dlc=0 dwc=0 vfbcv=-0.720472 noff=1 voffcv=0 acde=0.5 moin=15 wln=1 wl=0 wwn=1 ww=0 wwl=0 lln=1 ll=0 lwn=1 lw=0 lwl=0 llc=0 lwc=0 lwlc=0 wlc=0 wwc=0 wwlc=0 alpha0=0 alpha1=0 beta0=30 af=1.09369 kf=4.13676e-023 rsh=4 js=0.0001 jsw=0 
+ cj=0.00121101 mj=0.398913 pb=0.786344 cjsw=5.3952e-011 mjsw=2 tref=27 prt=0.628378 ute=-1.29285 kt1=-0.227499 kt1l=0 kt2=-0.0211773 ua1=5.21908e-010 ub1=9.72591e-019 uc1=2.64618e-011 at=10798.4 xti=3 tcj=0.00092022 tcjsw=-0.0079958 tpb=0.0022292 
+ tpbsw=-0.0087143 elm=5 xl=0 xw=0 ldif=1e-007 hdif=2.7e-007 lmlt=1 wmlt=1 rd=0 rdc=0 rs=0 rsc=0 php=0.8 cjgate=2e-014 n=1 

.model nmos_tkt2.12 nmos level=49 wmax=1e-005 wmin=1e-006 lmax=5e-007 lmin=3e-007 acm=2 version=3.2 mobmod=1 capmod=1 nqsmod=0 binunit=2 binflag=1 tox=5.05e-009 toxm=5.05e-009 xj=1e-007 nch=2.37707e+017 vth0=0.450123 lvth0=2.79026e-008 
+ wvth0=3.09035e-009 pvth0=-6.26889e-015 vfb=-0.62832 k1=0.392732 lk1=6.17893e-008 wk1=-1.00958e-007 pk1=2.61339e-014 k2=0.0514787 lk2=-3.94337e-008 wk2=2.76023e-009 pk2=-3.01426e-015 k3=0 k3b=0 w0=0 nlx=0 dvt0w=0 dvt1w=0 dvt2w=0 dvt0=0 dvt1=0 
+ dvt2=0 u0=0.0298893 lu0=3.53959e-009 wu0=-2.51919e-009 pu0=-1.93545e-015 ua=-5.05e-010 ub=1.73896e-018 lub=5.40078e-025 wub=-4.27624e-025 pub=-1.00393e-031 uc=1.14528e-010 luc=3.70879e-017 wuc=-7.66976e-017 puc=1.29249e-024 vsat=143933 
+ lvsat=-0.0187264 wvsat=-0.0180124 pvsat=3.77404e-009 a0=1.30902 la0=-3.64204e-007 wa0=2.5697e-007 pa0=-1.19674e-013 ags=-0.080968 lags=2.89592e-008 wags=7.49037e-008 pags=-2.22032e-014 b0=0 b1=0 keta=-0.00622539 lketa=-4.96004e-010 
+ wketa=1.44915e-008 pketa=-4.22619e-015 a1=0 a2=0.99 rdsw=10 prwg=0.2 prwb=-0.3 wr=1 wint=0 lint=0 dwg=0 dwb=0 voff=-0.100428 lvoff=3.05307e-009 wvoff=-7.31461e-008 pvoff=1.92282e-014 nfactor=0.377992 lnfactor=1.50492e-007 wnfactor=-5.12514e-007 
+ pnfactor=-8.32304e-014 eta0=-0.00484619 leta0=2.58813e-009 weta0=2.8926e-009 peta0=-4.84211e-016 etab=0.00206613 letab=-1.36177e-009 wetab=-7.71954e-010 petab=3.6195e-016 pclm=-0.0123225 lpclm=3.84886e-007 wpclm=8.17397e-007 ppclm=-3.23169e-013 
+ pdiblc1=0 pdiblc2=0.0196507 lpdiblc2=1.46329e-009 wpdiblc2=-6.35348e-009 ppdiblc2=-6.89866e-016 pdiblcb=-0.116243 lpdiblcb=4.14554e-008 wpdiblcb=2.05962e-007 ppdiblcb=-5.39871e-014 drout=0 pscbe1=7.70752e+008 pscbe2=1e-020 pvag=1.71485 
+ lpvag=-3.38253e-007 wpvag=-7.74811e-008 ppvag=-1.52956e-013 delta=0.01 ngate=1e+030 dsub=0 cit=0.00104355 lcit=-2.29622e-010 wcit=6.14629e-010 pcit=1.36209e-016 cdsc=0 cdscd=0 cdscb=0 xpart=0 cgso=3.15e-010 cgdo=3.15e-010 cgbo=1e-013 cgsl=0 cgdl=0 
+ ckappa=0.6 cf=0 clc=1e-007 cle=0.6 dlc=0 dwc=0 vfbcv=-0.720472 noff=1 voffcv=0 acde=0.5 moin=15 wln=1 wl=0 wwn=1 ww=0 wwl=0 lln=1 ll=0 lwn=1 lw=0 lwl=0 llc=0 lwc=0 lwlc=0 wlc=0 wwc=0 wwlc=0 alpha0=0 alpha1=0 beta0=30 af=1.09369 kf=4.13676e-023 
+ rsh=4 js=0.0001 jsw=0 cj=0.00121101 mj=0.398913 pb=0.786344 cjsw=5.3952e-011 mjsw=2 tref=27 prt=0.628378 ute=-1.29285 kt1=-0.227499 kt1l=0 kt2=-0.0211773 ua1=5.21908e-010 ub1=9.72591e-019 uc1=2.64618e-011 at=10798.4 xti=3 tcj=0.00092022 
+ tcjsw=-0.0079958 tpb=0.0022292 tpbsw=-0.0087143 elm=5 xl=0 xw=0 ldif=1e-007 hdif=2.7e-007 lmlt=1 wmlt=1 rd=0 rdc=0 rs=0 rsc=0 php=0.8 cjgate=2e-014 n=1 

.model nmos_tkt2.13 nmos level=49 wmax=1e-005 wmin=1e-006 lmax=1e-006 lmin=5e-007 acm=2 version=3.2 mobmod=1 capmod=1 nqsmod=0 binunit=2 binflag=1 tox=5.05e-009 toxm=5.05e-009 xj=1e-007 nch=2.37707e+017 vth0=0.44406 lvth0=3.09342e-008 
+ wvth0=-2.94917e-008 pvth0=1.00221e-014 vfb=-0.62832 k1=0.433003 lk1=4.1654e-008 wk1=-7.51611e-008 pk1=1.32355e-014 k2=-0.000891328 lk2=-1.32486e-008 wk2=1.64677e-008 pk2=-9.86801e-015 k3=0 k3b=0 w0=0 nlx=0 dvt0w=0 dvt1w=0 dvt2w=0 dvt0=0 dvt1=0 
+ dvt2=0 u0=0.0331092 lu0=1.92966e-009 wu0=-6.52586e-009 pu0=6.7888e-017 ua=-5.05e-010 ub=1.57658e-018 lub=6.21268e-025 wub=-1.34006e-025 pub=-2.47202e-031 uc=1.05824e-011 luc=8.90608e-017 wuc=-4.28538e-018 puc=-3.49136e-023 vsat=893520 
+ lvsat=-0.39352 wvsat=0.0104643 pvsat=-1.04643e-008 a0=1.78158 la0=-6.00483e-007 wa0=-7.29115e-008 pa0=4.52668e-014 ags=-0.0169503 lags=-3.04973e-009 wags=-3.04972e-008 pags=3.04972e-014 b0=0 b1=0 keta=0.0251191 lketa=-1.61682e-008 
+ wketa=-5.823e-009 pketa=5.93107e-015 a1=0 a2=0.99 rdsw=10 prwg=0.2 prwb=-0.3 wr=1 wint=0 lint=0 dwg=0 dwb=0 voff=-0.104122 lvoff=4.90012e-009 wvoff=-2.92025e-008 pvoff=-2.74362e-015 nfactor=0.34686 lnfactor=1.66058e-007 wnfactor=-3.4686e-007 
+ pnfactor=-1.66058e-013 eta0=0.00201148 leta0=-8.40701e-010 weta0=-3.3811e-009 peta0=2.65264e-015 etab=8.286e-005 letab=-3.7014e-010 wetab=3.78002e-010 petab=-2.13028e-016 pclm=-1.84634 lpclm=1.3019e-006 wpclm=1.09178e-005 ppclm=-5.37339e-012 
+ pdiblc1=0 pdiblc2=0.0455599 lpdiblc2=-1.14913e-008 wpdiblc2=1.39596e-007 ppdiblc2=-7.36646e-014 pdiblcb=0.401248 lpdiblcb=-2.1729e-007 wpdiblcb=-6.59041e-008 ppdiblcb=8.19461e-014 drout=0 pscbe1=7.70752e+008 pscbe2=1e-020 pvag=1.18388 
+ lpvag=-7.27718e-008 wpvag=-1.83883e-006 ppvag=7.27718e-013 delta=0.01 ngate=1e+030 dsub=0 cit=0.00114572 lcit=-2.80708e-010 wcit=-1.0372e-009 pcit=9.62122e-016 cdsc=0 cdscd=-8.43816e-006 lcdscd=4.21908e-012 wcdscd=8.43815e-011 pcdscd=-4.21908e-017 
+ cdscb=0 xpart=0 cgso=3.15e-010 cgdo=3.15e-010 cgbo=1e-013 cgsl=0 cgdl=0 ckappa=0.6 cf=0 clc=1e-007 cle=0.6 dlc=0 dwc=0 vfbcv=-0.720472 noff=1 voffcv=0 acde=0.5 moin=15 wln=1 wl=0 wwn=1 ww=0 wwl=0 lln=1 ll=0 lwn=1 lw=0 lwl=0 llc=0 lwc=0 lwlc=0 
+ wlc=0 wwc=0 wwlc=0 alpha0=0 alpha1=0 beta0=30 af=1.09369 kf=4.13676e-023 rsh=4 js=0.0001 jsw=0 cj=0.00121101 mj=0.398913 pb=0.786344 cjsw=5.3952e-011 mjsw=2 tref=27 prt=0.628378 ute=-1.29285 kt1=-0.227499 kt1l=0 kt2=-0.0211773 ua1=5.21908e-010 
+ ub1=9.72591e-019 uc1=2.64618e-011 at=10798.4 xti=3 tcj=0.00092022 tcjsw=-0.0079958 tpb=0.0022292 tpbsw=-0.0087143 elm=5 xl=0 xw=0 ldif=1e-007 hdif=2.7e-007 lmlt=1 wmlt=1 rd=0 rdc=0 rs=0 rsc=0 php=0.8 cjgate=2e-014 n=1 

.model nmos_tkt2.14 nmos level=49 wmax=1e-005 wmin=1e-006 lmax=1e-005 lmin=1e-006 acm=2 version=3.2 mobmod=1 capmod=1 nqsmod=0 binunit=2 binflag=1 tox=5.05e-009 toxm=5.05e-009 xj=1e-007 nch=2.37707e+017 vth0=0.393012 lvth0=8.19817e-008 
+ wvth0=-7.54267e-009 pvth0=-1.19269e-014 vfb=-0.62832 k1=0.438402 lk1=3.62546e-008 wk1=-1.82624e-008 pk1=-4.36632e-014 k2=0.00485961 lk2=-1.89995e-008 wk2=-5.26599e-009 pk2=1.18657e-014 k3=0 k3b=0 w0=0 nlx=0 dvt0w=0 dvt1w=0 dvt2w=0 dvt0=0 dvt1=0 
+ dvt2=0 u0=0.0338295 lu0=1.20932e-009 wu0=-6.68252e-009 pu0=2.24542e-016 ua=-5.05003e-010 wua=3.02227e-020 pua=-3.02227e-026 ub=1.73125e-018 lub=4.66596e-025 wub=-1.86369e-025 pub=-1.94838e-031 uc=3.56312e-011 luc=6.4012e-017 wuc=-1.73979e-017 
+ puc=-2.18011e-023 vsat=500000 a0=0.439942 la0=7.41153e-007 wa0=7.28672e-008 pa0=-1.00512e-013 ags=0.0244444 lags=-4.44444e-008 b0=0 b1=0 keta=0.00905137 lketa=-1.00541e-010 wketa=1.69601e-009 pketa=-1.58794e-015 a1=0 a2=0.99 rdsw=10 prwg=0.2 
+ prwb=-0.3 wr=1 wint=0 lint=0 dwg=0 dwb=0 voff=-0.0957097 lvoff=-3.51197e-009 wvoff=-3.99204e-008 pvoff=7.9743e-015 nfactor=0.394516 lnfactor=1.18402e-007 wnfactor=-3.94516e-007 pnfactor=-1.18402e-013 eta0=-0.000135788 leta0=1.30656e-009 
+ weta0=4.77767e-010 peta0=-1.20623e-015 etab=3.192e-005 letab=-3.192e-010 wetab=-1.83304e-011 petab=1.83304e-016 pclm=5.61605 pdiblc1=0 pdiblc2=0.107326 lpdiblc2=-7.32572e-008 wpdiblc2=-7.32572e-009 ppdiblc2=7.32572e-014 pdiblcb=0.201783 
+ lpdiblcb=-1.78245e-008 wpdiblcb=-1.78245e-009 ppdiblcb=1.78245e-014 drout=0 pscbe1=7.70752e+008 pscbe2=1e-020 pvag=-0.123457 lpvag=1.23457e-006 wpvag=1.23457e-007 ppvag=-1.23457e-012 delta=0.01 ngate=1e+030 dsub=0 cit=0.000795005 lcit=7.00108e-011 
+ wcit=2.01504e-010 pcit=-2.7658e-016 cdsc=0 cdscd=4.23738e-005 lcdscd=-4.65929e-011 wcdscd=-4.65929e-011 pcdscd=8.87837e-017 cdscb=0 xpart=0 cgso=3.15e-010 cgdo=3.15e-010 cgbo=1e-013 cgsl=0 cgdl=0 ckappa=0.6 cf=0 clc=1e-007 cle=0.6 dlc=0 dwc=0 
+ vfbcv=-0.720472 noff=1 voffcv=0 acde=0.5 moin=15 wln=1 wl=0 wwn=1 ww=0 wwl=0 lln=1 ll=0 lwn=1 lw=0 lwl=0 llc=0 lwc=0 lwlc=0 wlc=0 wwc=0 wwlc=0 alpha0=0 alpha1=0 beta0=30 af=1.09369 kf=4.13676e-023 rsh=4 js=0.0001 jsw=0 cj=0.00121101 mj=0.398913 
+ pb=0.786344 cjsw=5.3952e-011 mjsw=2 tref=27 prt=0.628378 ute=-1.29285 kt1=-0.227499 kt1l=0 kt2=-0.0211773 ua1=5.21908e-010 ub1=9.72591e-019 uc1=2.64618e-011 at=10798.4 xti=3 tcj=0.00092022 tcjsw=-0.0079958 tpb=0.0022292 tpbsw=-0.0087143 elm=5 xl=0 
+ xw=0 ldif=1e-007 hdif=2.7e-007 lmlt=1 wmlt=1 rd=0 rdc=0 rs=0 rsc=0 php=0.8 cjgate=2e-014 n=1 

.model nmos_tkt2.15 nmos level=49 wmax=1e-005 wmin=1e-006 lmax=2e-005 lmin=1e-005 acm=2 version=3.2 mobmod=1 capmod=1 nqsmod=0 binunit=2 binflag=1 tox=5.05e-009 toxm=5.05e-009 xj=1e-007 nch=2.37707e+017 vth0=0.401211 wvth0=-8.73536e-009 vfb=-0.62832 
+ k1=0.442028 wk1=-2.26287e-008 k2=0.00295966 wk2=-4.07942e-009 k3=0 k3b=0 w0=0 nlx=0 dvt0w=0 dvt1w=0 dvt2w=0 dvt0=0 dvt1=0 dvt2=0 u0=0.0339504 wu0=-6.66006e-009 ua=-5.05003e-010 wua=2.72005e-020 ub=1.77791e-018 wub=-2.05853e-025 uc=4.20324e-011 
+ wuc=-1.9578e-017 vsat=500000 a0=0.514057 wa0=6.2816e-008 ags=0.02 b0=0 b1=0 keta=0.00904131 wketa=1.53722e-009 a1=0 a2=0.99 rdsw=10 prwg=0.2 prwb=-0.3 wr=1 wint=0 lint=0 dwg=0 dwb=0 voff=-0.0960609 wvoff=-3.9123e-008 nfactor=0.406356 
+ wnfactor=-4.06356e-007 eta0=-5.13133e-006 weta0=3.57144e-010 etab=0 pclm=5 pdiblc1=0 pdiblc2=0.1 pdiblcb=0.2 drout=0 pscbe1=7.70752e+008 pscbe2=1e-020 pvag=0 delta=0.01 ngate=1e+030 dsub=0 cit=0.000802006 wcit=1.73846e-010 cdsc=0 
+ cdscd=3.77145e-005 wcdscd=-3.77145e-011 cdscb=0 xpart=0 cgso=3.15e-010 cgdo=3.15e-010 cgbo=1e-013 cgsl=0 cgdl=0 ckappa=0.6 cf=0 clc=1e-007 cle=0.6 dlc=0 dwc=0 vfbcv=-0.720472 noff=1 voffcv=0 acde=0.5 moin=15 wln=1 wl=0 wwn=1 ww=0 wwl=0 lln=1 ll=0 
+ lwn=1 lw=0 lwl=0 llc=0 lwc=0 lwlc=0 wlc=0 wwc=0 wwlc=0 alpha0=0 alpha1=0 beta0=30 af=1.09369 kf=4.13676e-023 rsh=4 js=0.0001 jsw=0 cj=0.00121101 mj=0.398913 pb=0.786344 cjsw=5.3952e-011 mjsw=2 tref=27 prt=0.628378 ute=-1.29285 kt1=-0.227499 kt1l=0 
+ kt2=-0.0211773 ua1=5.21908e-010 ub1=9.72591e-019 uc1=2.64618e-011 at=10798.4 xti=3 tcj=0.00092022 tcjsw=-0.0079958 tpb=0.0022292 tpbsw=-0.0087143 elm=5 xl=0 xw=0 ldif=1e-007 hdif=2.7e-007 lmlt=1 wmlt=1 rd=0 rdc=0 rs=0 rsc=0 php=0.8 cjgate=2e-014 
+ n=1 

.model nmos_tkt2.16 nmos level=49 wmax=0.0001 wmin=1e-005 lmax=3e-007 lmin=2.4e-007 acm=2 version=3.2 mobmod=1 capmod=1 nqsmod=0 binunit=2 binflag=1 tox=5.05e-009 toxm=5.05e-009 xj=1e-007 nch=2.37707e+017 vth0=0.524838 lvth0=4.954e-009 vfb=-0.62832 
+ k1=0.740441 lk1=-4.29386e-008 k2=-0.0221721 lk2=-1.7557e-008 k3=0 k3b=0 w0=0 nlx=0 dvt0w=0 dvt1w=0 dvt2w=0 dvt0=0 dvt1=0 dvt2=0 u0=-0.0650768 lu0=3.17603e-008 ua=-9.2017e-009 lua=2.60901e-015 ub=-8.28378e-020 lub=1.06375e-024 uc=-4.54576e-010 
+ luc=2.05648e-016 vsat=86491.9 lvsat=-0.00165703 a0=0.608001 la0=-1.58157e-007 ags=0.0867536 lags=-2.13305e-008 b0=0 b1=0 keta=-0.0275982 lketa=5.92795e-009 a1=0 a2=0.99 rdsw=10 prwg=1.8 lprwg=-4.8e-007 prwb=-2.7 lprwb=7.2e-007 wr=1 wint=0 lint=0 
+ dwg=0 dwb=0 voff=-0.0535113 lvoff=-1.12934e-008 nfactor=2.70474 lnfactor=-5.71232e-007 eta0=-0.0151263 leta0=5.71051e-009 etab=0.00123707 letab=-1.10002e-009 pclm=0.588398 lpclm=1.96875e-007 pdiblc1=0 pdiblc2=0.00780621 lpdiblc2=4.75704e-009 
+ pdiblcb=-0.310717 lpdiblcb=1.00578e-007 drout=0 pscbe1=7.70752e+008 pscbe2=1e-020 pvag=0.357791 lpvag=5.12431e-008 delta=0.01 ngate=1e+030 dsub=0 cit=-0.00289387 lcit=9.83664e-010 cdsc=0 cdscd=-0.000164846 lcdscd=4.94539e-011 cdscb=0 xpart=0 
+ cgso=3.15e-010 cgdo=3.15e-010 cgbo=1e-013 cgsl=0 cgdl=0 ckappa=0.6 cf=0 clc=1e-007 cle=0.6 dlc=0 dwc=0 vfbcv=-0.720472 noff=1 voffcv=0 acde=0.5 moin=15 wln=1 wl=0 wwn=1 ww=0 wwl=0 lln=1 ll=0 lwn=1 lw=0 lwl=0 llc=0 lwc=0 lwlc=0 wlc=0 wwc=0 wwlc=0 
+ alpha0=0 alpha1=0 beta0=30 af=1.09369 kf=4.13676e-023 rsh=4 js=0.0001 jsw=0 cj=0.00121101 mj=0.398913 pb=0.786344 cjsw=5.3952e-011 mjsw=2 tref=27 prt=0.628378 ute=-1.29285 kt1=-0.227499 kt1l=0 kt2=-0.0211773 ua1=5.21908e-010 ub1=9.72591e-019 
+ uc1=2.64618e-011 at=10798.4 xti=3 tcj=0.00092022 tcjsw=-0.0079958 tpb=0.0022292 tpbsw=-0.0087143 elm=5 xl=0 xw=0 ldif=1e-007 hdif=2.7e-007 lmlt=1 wmlt=1 rd=0 rdc=0 rs=0 rsc=0 php=0.8 cjgate=2e-014 n=1 

.model nmos_tkt2.17 nmos level=49 wmax=0.0001 wmin=1e-005 lmax=5e-007 lmin=3e-007 acm=2 version=3.2 mobmod=1 capmod=1 nqsmod=0 binunit=2 binflag=1 tox=5.05e-009 toxm=5.05e-009 xj=1e-007 nch=2.37707e+017 vth0=0.450432 lvth0=2.72757e-008 vfb=-0.62832 
+ k1=0.382636 lk1=6.44027e-008 k2=0.0517548 lk2=-3.97351e-008 k3=0 k3b=0 w0=0 nlx=0 dvt0w=0 dvt1w=0 dvt2w=0 dvt0=0 dvt1=0 dvt2=0 u0=0.0296374 lu0=3.34605e-009 ua=-5.05e-010 ub=1.6962e-018 lub=5.30038e-025 uc=1.06858e-010 luc=3.72171e-017 vsat=142132 
+ lvsat=-0.018349 a0=1.33472 la0=-3.76172e-007 ags=-0.0734777 lags=2.67388e-008 b0=0 b1=0 keta=-0.00477624 lketa=-9.18622e-010 a1=0 a2=0.99 rdsw=10 prwg=0.2 prwb=-0.3 wr=1 wint=0 lint=0 dwg=0 dwb=0 voff=-0.107742 lvoff=4.97589e-009 nfactor=0.32674 
+ lnfactor=1.42169e-007 eta0=-0.00455692 leta0=2.53971e-009 etab=0.00198893 letab=-1.32558e-009 pclm=0.0694172 lpclm=3.5257e-007 pdiblc1=0 pdiblc2=0.0190153 lpdiblc2=1.39431e-009 pdiblcb=-0.0956465 lpdiblcb=3.60566e-008 drout=0 pscbe1=7.70752e+008 
+ pscbe2=1e-020 pvag=1.7071 lpvag=-3.53549e-007 delta=0.01 ngate=1e+030 dsub=0 cit=0.00110501 lcit=-2.16001e-010 cdsc=0 cdscd=0 cdscb=0 xpart=0 cgso=3.15e-010 cgdo=3.15e-010 cgbo=1e-013 cgsl=0 cgdl=0 ckappa=0.6 cf=0 clc=1e-007 cle=0.6 dlc=0 dwc=0 
+ vfbcv=-0.720472 noff=1 voffcv=0 acde=0.5 moin=15 wln=1 wl=0 wwn=1 ww=0 wwl=0 lln=1 ll=0 lwn=1 lw=0 lwl=0 llc=0 lwc=0 lwlc=0 wlc=0 wwc=0 wwlc=0 alpha0=0 alpha1=0 beta0=30 af=1.09369 kf=4.13676e-023 rsh=4 js=0.0001 jsw=0 cj=0.00121101 mj=0.398913 
+ pb=0.786344 cjsw=5.3952e-011 mjsw=2 tref=27 prt=0.628378 ute=-1.29285 kt1=-0.227499 kt1l=0 kt2=-0.0211773 ua1=5.21908e-010 ub1=9.72591e-019 uc1=2.64618e-011 at=10798.4 xti=3 tcj=0.00092022 tcjsw=-0.0079958 tpb=0.0022292 tpbsw=-0.0087143 elm=5 xl=0 
+ xw=0 ldif=1e-007 hdif=2.7e-007 lmlt=1 wmlt=1 rd=0 rdc=0 rs=0 rsc=0 php=0.8 cjgate=2e-014 n=1 

.model nmos_tkt2.18 nmos level=49 wmax=0.0001 wmin=1e-005 lmax=1e-006 lmin=5e-007 acm=2 version=3.2 mobmod=1 capmod=1 nqsmod=0 binunit=2 binflag=1 tox=5.05e-009 toxm=5.05e-009 xj=1e-007 nch=2.37707e+017 vth0=0.441111 vfb=-0.62832 k1=0.425487 
+ lk1=4.29775e-008 k2=0.000755444 lk2=-1.42354e-008 k3=0 k3b=0 w0=0 nlx=0 dvt0w=0 dvt1w=0 dvt2w=0 dvt0=0 dvt1=0 dvt2=0 u0=0.0324566 lu0=1.93645e-009 ua=-5.05e-010 ub=1.56318e-018 lub=5.96548e-025 uc=1.01539e-011 luc=8.55694e-017 vsat=894566 
+ lvsat=-0.394566 a0=1.77429 la0=-5.95956e-007 ags=-0.02 b0=0 b1=0 keta=0.0245368 lketa=-1.55751e-008 a1=0 a2=0.99 rdsw=10 prwg=0.2 prwb=-0.3 wr=1 wint=0 lint=0 dwg=0 dwb=0 voff=-0.107042 lvoff=4.62575e-009 nfactor=0.312174 lnfactor=1.49452e-007 
+ eta0=0.00167337 leta0=-5.75438e-010 etab=0.00012066 letab=-3.91443e-010 pclm=-0.754556 lpclm=7.64556e-007 pdiblc1=0 pdiblc2=0.0595195 lpdiblc2=-1.88578e-008 pdiblcb=0.394658 lpdiblcb=-2.09095e-007 drout=0 pscbe1=7.70752e+008 pscbe2=1e-020 pvag=1 
+ delta=0.01 ngate=1e+030 dsub=0 cit=0.001042 lcit=-1.84496e-010 cdsc=0 cdscd=0 cdscb=0 xpart=0 cgso=3.15e-010 cgdo=3.15e-010 cgbo=1e-013 cgsl=0 cgdl=0 ckappa=0.6 cf=0 clc=1e-007 cle=0.6 dlc=0 dwc=0 vfbcv=-0.720472 noff=1 voffcv=0 acde=0.5 moin=15 
+ wln=1 wl=0 wwn=1 ww=0 wwl=0 lln=1 ll=0 lwn=1 lw=0 lwl=0 llc=0 lwc=0 lwlc=0 wlc=0 wwc=0 wwlc=0 alpha0=0 alpha1=0 beta0=30 af=1.09369 kf=4.13676e-023 rsh=4 js=0.0001 jsw=0 cj=0.00121101 mj=0.398913 pb=0.786344 cjsw=5.3952e-011 mjsw=2 tref=27 
+ prt=0.628378 ute=-1.29285 kt1=-0.227499 kt1l=0 kt2=-0.0211773 ua1=5.21908e-010 ub1=9.72591e-019 uc1=2.64618e-011 at=10798.4 xti=3 tcj=0.00092022 tcjsw=-0.0079958 tpb=0.0022292 tpbsw=-0.0087143 elm=5 xl=0 xw=0 ldif=1e-007 hdif=2.7e-007 lmlt=1 
+ wmlt=1 rd=0 rdc=0 rs=0 rsc=0 php=0.8 cjgate=2e-014 n=1 

.model nmos_tkt2.19 nmos level=49 wmax=0.0001 wmin=1e-005 lmax=1e-005 lmin=1e-006 acm=2 version=3.2 mobmod=1 capmod=1 nqsmod=0 binunit=2 binflag=1 tox=5.05e-009 toxm=5.05e-009 xj=1e-007 nch=2.37707e+017 vth0=0.392258 lvth0=8.0789e-008 vfb=-0.62832 
+ k1=0.436576 lk1=3.18883e-008 k2=0.00433301 lk2=-1.7813e-008 k3=0 k3b=0 w0=0 nlx=0 dvt0w=0 dvt1w=0 dvt2w=0 dvt0=0 dvt1=0 dvt2=0 u0=0.0331613 lu0=1.23178e-009 ua=-5.05e-010 ub=1.71261e-018 lub=4.47112e-025 uc=3.38914e-011 luc=6.18319e-017 
+ vsat=500000 a0=0.447229 la0=7.31102e-007 ags=0.0244444 lags=-4.44444e-008 b0=0 b1=0 keta=0.00922097 lketa=-2.59335e-010 a1=0 a2=0.99 rdsw=10 prwg=0.2 prwb=-0.3 wr=1 wint=0 lint=0 dwg=0 dwb=0 voff=-0.0997018 lvoff=-2.71454e-009 nfactor=0.355064 
+ lnfactor=1.06562e-007 eta0=-8.80112e-005 leta0=1.18594e-009 etab=3.0087e-005 letab=-3.00869e-010 pclm=5.55445 pdiblc1=0 pdiblc2=0.106593 lpdiblc2=-6.59314e-008 pdiblcb=0.201604 lpdiblcb=-1.6042e-008 drout=0 pscbe1=7.70752e+008 pscbe2=1e-020 
+ pvag=-0.111111 lpvag=1.11111e-006 delta=0.01 ngate=1e+030 dsub=0 cit=0.000815155 lcit=4.23528e-011 cdsc=0 cdscd=3.77145e-005 lcdscd=-3.77145e-011 cdscb=0 xpart=0 cgso=3.15e-010 cgdo=3.15e-010 cgbo=1e-013 cgsl=0 cgdl=0 ckappa=0.6 cf=0 clc=1e-007 
+ cle=0.6 dlc=0 dwc=0 vfbcv=-0.720472 noff=1 voffcv=0 acde=0.5 moin=15 wln=1 wl=0 wwn=1 ww=0 wwl=0 lln=1 ll=0 lwn=1 lw=0 lwl=0 llc=0 lwc=0 lwlc=0 wlc=0 wwc=0 wwlc=0 alpha0=0 alpha1=0 beta0=30 af=1.09369 kf=4.13676e-023 rsh=4 js=0.0001 jsw=0 
+ cj=0.00121101 mj=0.398913 pb=0.786344 cjsw=5.3952e-011 mjsw=2 tref=27 prt=0.628378 ute=-1.29285 kt1=-0.227499 kt1l=0 kt2=-0.0211773 ua1=5.21908e-010 ub1=9.72591e-019 uc1=2.64618e-011 at=10798.4 xti=3 tcj=0.00092022 tcjsw=-0.0079958 tpb=0.0022292 
+ tpbsw=-0.0087143 elm=5 xl=0 xw=0 ldif=1e-007 hdif=2.7e-007 lmlt=1 wmlt=1 rd=0 rdc=0 rs=0 rsc=0 php=0.8 cjgate=2e-014 n=1 

.model nmos_tkt2.20 nmos level=49 wmax=0.0001 wmin=1e-005 lmax=2e-005 lmin=1e-005 acm=2 version=3.2 mobmod=1 capmod=1 nqsmod=0 binunit=2 binflag=1 tox=5.05e-009 toxm=5.05e-009 xj=1e-007 nch=2.37707e+017 vth0=0.400337 vfb=-0.62832 k1=0.439765 
+ k2=0.00255171 k3=0 k3b=0 w0=0 nlx=0 dvt0w=0 dvt1w=0 dvt2w=0 dvt0=0 dvt1=0 dvt2=0 u0=0.0332844 ua=-5.05e-010 ub=1.75732e-018 uc=4.00746e-011 vsat=500000 a0=0.520339 ags=0.02 b0=0 b1=0 keta=0.00919504 a1=0 a2=0.99 rdsw=10 prwg=0.2 prwb=-0.3 wr=1 
+ wint=0 lint=0 dwg=0 dwb=0 voff=-0.0999732 nfactor=0.36572 eta0=3.05831e-005 etab=0 pclm=5 pdiblc1=0 pdiblc2=0.1 pdiblcb=0.2 drout=0 pscbe1=7.70752e+008 pscbe2=1e-020 pvag=0 delta=0.01 ngate=1e+030 dsub=0 cit=0.000819391 cdsc=0 cdscd=3.39431e-005 
+ cdscb=0 xpart=0 cgso=3.15e-010 cgdo=3.15e-010 cgbo=1e-013 cgsl=0 cgdl=0 ckappa=0.6 cf=0 clc=1e-007 cle=0.6 dlc=0 dwc=0 vfbcv=-0.720472 noff=1 voffcv=0 acde=0.5 moin=15 wln=1 wl=0 wwn=1 ww=0 wwl=0 lln=1 ll=0 lwn=1 lw=0 lwl=0 llc=0 lwc=0 lwlc=0 
+ wlc=0 wwc=0 wwlc=0 alpha0=0 alpha1=0 beta0=30 af=1.09369 kf=4.13676e-023 rsh=4 js=0.0001 jsw=0 cj=0.00121101 mj=0.398913 pb=0.786344 cjsw=5.3952e-011 mjsw=2 tref=27 prt=0.628378 ute=-1.29285 kt1=-0.227499 kt1l=0 kt2=-0.0211773 ua1=5.21908e-010 
+ ub1=9.72591e-019 uc1=2.64618e-011 at=10798.4 xti=3 tcj=0.00092022 tcjsw=-0.0079958 tcjswg=0.0019057 tpb=0.0022292 tpbsw=-0.0087143 elm=5 xl=0 xw=0 ldif=1e-007 hdif=2.7e-007 lmlt=1 wmlt=1 rd=0 rdc=0 rs=0 rsc=0 php=0.8 cjgate=2e-014 n=1 

.model pmos_tkt2.1 pmos level=49 wmax=4e-007 wmin=3e-007 lmax=3e-007 lmin=2.4e-007 acm=2 version=3.2 mobmod=1 capmod=1 nqsmod=0 binunit=2 binflag=1 tox=5.05e-009 toxm=5.05e-009 xj=1e-007 nch=3.29929e+017 vth0=0.65295 lvth0=-3.05316e-007 
+ wvth0=-3.19176e-007 pvth0=9.26828e-014 vfb=-0.62832 k1=-16.3926 lk1=4.06555e-006 wk1=6.72786e-006 pk1=-1.62616e-012 k2=6.02375 lk2=-1.45763e-006 wk2=-2.40895e-006 pk2=5.78483e-013 k3=0 k3b=0 w0=0 nlx=0 dvt0w=0 dvt1w=0 dvt2w=0 dvt0=0 dvt1=0 dvt2=0 
+ u0=-0.0123383 lu0=6.79714e-009 wu0=5.12668e-009 pu0=-1.91716e-015 ua=-5.48157e-009 lua=1.92345e-015 wua=1.28527e-015 pua=-4.68576e-022 ub=1.86134e-018 lub=1.74302e-025 wub=-4.87069e-025 pub=1.59584e-032 uc=6.17421e-011 luc=3.86294e-017 
+ wuc=-8.61046e-017 puc=4.5408e-024 vsat=2.10867e+006 lvsat=-0.365553 wvsat=-0.5331 pvsat=9.68291e-008 a0=20.8585 la0=-5.20046e-006 wa0=-7.65967e-006 pa0=2.00295e-012 ags=0.296226 lags=-6.48678e-008 wags=-1.1049e-007 pags=2.59471e-014 b0=0 b1=0 
+ keta=0.514471 lketa=-1.35843e-007 wketa=-1.88787e-007 pketa=5.04709e-014 a1=0 a2=0.4 rdsw=10 prwg=0.2 prwb=-0.3 wr=1 wint=0 lint=0 dwg=0 dwb=0 voff=-0.156381 lvoff=-9.44537e-009 wvoff=5.62913e-008 pvoff=-6.75084e-015 nfactor=39.7845 
+ lnfactor=-1.09185e-005 wnfactor=-1.31577e-005 pnfactor=3.70595e-012 eta0=0.0982337 leta0=-2.45495e-008 weta0=-4.09287e-008 peta0=1.08024e-014 etab=-0.0244062 letab=5.55831e-009 wetab=9.36095e-009 petab=-2.29141e-015 pclm=54.0191 
+ lpclm=-1.23141e-005 wpclm=-1.4905e-005 ppclm=3.51485e-012 pdiblc1=0 pdiblc2=-0.80113 lpdiblc2=1.96373e-007 wpdiblc2=3.13624e-007 ppdiblc2=-7.64995e-014 pdiblcb=12.5938 lpdiblcb=-3.35836e-006 wpdiblcb=-4.31789e-006 ppdiblcb=1.15144e-012 drout=0 
+ pscbe1=7.70752e+008 pscbe2=1e-020 pvag=-19 lpvag=4.8e-006 wpvag=6e-006 ppvag=-1.44e-012 delta=0.01 ngate=1e+030 dsub=0 cit=-0.00502783 lcit=2.89689e-009 wcit=-7.40658e-010 pcit=-3.67077e-016 cdsc=0 cdscd=-0.0043307 lcdscd=1.06137e-009 
+ wcdscd=1.7606e-009 pcdscd=-4.28252e-016 cdscb=0 xpart=0 cgso=2.2653e-010 cgdo=2.2653e-010 cgbo=1e-013 cgsl=0 cgdl=0 ckappa=0.6 cf=0 clc=1e-007 cle=0.6 dlc=0 dwc=0 vfbcv=-0.826159 noff=1 voffcv=0 acde=0.5 moin=15 wln=1 wl=0 wwn=1 ww=0 wwl=0 lln=1 
+ ll=0 lwn=1 lw=0 lwl=0 llc=0 lwc=0 lwlc=0 wlc=0 wwc=0 wwlc=0 alpha0=0 alpha1=0 beta0=30 af=1.1021 kf=1.74179e-023 rsh=3 js=0.0001 jsw=0 cj=0.00150656 mj=0.403022 pb=0.790743 cjsw=1.18641e-010 mjsw=2 tref=27 prt=-149.998 ute=-0.950103 kt1=-0.257006 
+ kt1l=0 kt2=-0.0222175 ua1=1.29549e-010 ub1=-1.58953e-018 uc1=-4.01361e-011 at=-50000 xti=3 tcj=0.00075544 tcjsw=0.0017757 tpb=0.0016635 tpbsw=-0.0013729 elm=5 xl=0 xw=0 ldif=1e-007 hdif=2.7e-007 lmlt=1 wmlt=1 rd=0 rdc=0 rs=0 rsc=0 php=0.8 
+ cjgate=2e-014 n=1 

.model pmos_tkt2.2 pmos level=49 wmax=4e-007 wmin=3e-007 lmax=5e-007 lmin=3e-007 acm=2 version=3.2 mobmod=1 capmod=1 nqsmod=0 binunit=2 binflag=1 tox=5.05e-009 toxm=5.05e-009 xj=1e-007 nch=3.29929e+017 vth0=-0.534034 lvth0=5.07794e-008 
+ wvth0=4.38008e-008 pvth0=-1.62103e-014 vfb=-0.62832 k1=5.489 lk1=-2.49892e-006 wk1=-2.01343e-006 pk1=9.96232e-013 k2=-1.74334 lk2=8.72499e-007 wk2=6.85196e-007 pk2=-3.49761e-013 k3=0 k3b=0 w0=0 nlx=0 dvt0w=0 dvt1w=0 dvt2w=0 dvt0=0 dvt1=0 dvt2=0 
+ u0=0.00451686 lu0=1.74059e-009 wu0=5.62278e-010 pu0=-5.47841e-016 ua=4.16255e-010 lua=1.54096e-016 wua=-4.61132e-017 pua=-6.91598e-023 ub=-1.83716e-018 lub=1.28385e-024 wub=5.83508e-025 pub=-3.05215e-031 uc=-4.10477e-010 luc=1.80295e-016 
+ wuc=1.00419e-016 puc=-5.14163e-023 vsat=-376325 lvsat=0.379945 wvsat=0.215514 pvsat=-1.27755e-007 a0=-3.6726 la0=2.15888e-006 wa0=1.52929e-006 pa0=-7.53733e-013 ags=-0.261643 lags=1.02493e-007 wags=9.26573e-008 pags=-3.49972e-014 b0=0 b1=0 
+ keta=-0.151562 lketa=6.39669e-008 wketa=5.28648e-008 pketa=-2.20247e-014 a1=0 a2=0.4 rdsw=10 prwg=0.2 prwb=-0.3 wr=1 wint=0 lint=0 dwg=0 dwb=0 voff=0.193433 lvoff=-1.1439e-007 wvoff=-1.33105e-007 pvoff=5.00682e-014 nfactor=-0.0840091 
+ lnfactor=1.042e-006 wnfactor=1.20677e-006 pnfactor=-6.03386e-013 eta0=-0.02101 leta0=1.12236e-008 weta0=7.17308e-009 peta0=-3.62811e-015 etab=0.00703988 letab=-3.87553e-009 wetab=-2.08331e-009 petab=1.14186e-015 pclm=-17.4756 lpclm=9.1343e-006 
+ wpclm=7.35275e-006 ppclm=-3.16248e-012 pdiblc1=0 pdiblc2=0.233168 lpdiblc2=-1.13917e-007 wpdiblc2=-9.1932e-008 ppdiblc2=4.51673e-014 pdiblcb=-1.59736 lpdiblcb=8.98975e-007 wpdiblcb=7.19063e-007 ppdiblcb=-3.59648e-013 drout=0 pscbe1=7.70752e+008 
+ pscbe2=1e-020 pvag=7 lpvag=-3e-006 wpvag=-1.8e-006 ppvag=9e-013 delta=0.01 ngate=1e+030 dsub=0 cit=-0.00600879 lcit=3.19118e-009 wcit=1.0266e-009 pcit=-8.97256e-016 cdsc=0 cdscd=0.00157033 lcdscd=-7.08935e-010 wcdscd=-6.13982e-010 
+ pcdscd=2.84122e-016 cdscb=0 xpart=0 cgso=2.2653e-010 cgdo=2.2653e-010 cgbo=1e-013 cgsl=0 cgdl=0 ckappa=0.6 cf=0 clc=1e-007 cle=0.6 dlc=0 dwc=0 vfbcv=-0.826159 noff=1 voffcv=0 acde=0.5 moin=15 wln=1 wl=0 wwn=1 ww=0 wwl=0 lln=1 ll=0 lwn=1 lw=0 lwl=0 
+ llc=0 lwc=0 lwlc=0 wlc=0 wwc=0 wwlc=0 alpha0=0 alpha1=0 beta0=30 af=1.1021 kf=1.74179e-023 rsh=3 js=0.0001 jsw=0 cj=0.00150656 mj=0.403022 pb=0.790743 cjsw=1.18641e-010 mjsw=2 tref=27 prt=-149.998 ute=-0.950103 kt1=-0.257006 kt1l=0 kt2=-0.0222175 
+ ua1=1.29549e-010 ub1=-1.58953e-018 uc1=-4.01361e-011 at=-50000 xti=3 tcj=0.00075544 tcjsw=0.0017757 tpb=0.0016635 tpbsw=-0.0013729 elm=5 xl=0 xw=0 ldif=1e-007 hdif=2.7e-007 lmlt=1 wmlt=1 rd=0 rdc=0 rs=0 rsc=0 php=0.8 cjgate=2e-014 n=1 

.model pmos_tkt2.3 pmos level=49 wmax=4e-007 wmin=3e-007 lmax=1e-006 lmin=5e-007 acm=2 version=3.2 mobmod=1 capmod=1 nqsmod=0 binunit=2 binflag=1 tox=5.05e-009 toxm=5.05e-009 xj=1e-007 nch=3.29929e+017 vth0=-0.674049 lvth0=1.20787e-007 
+ wvth0=8.94468e-008 pvth0=-3.90334e-014 vfb=-0.62832 k1=0.644477 lk1=-7.66585e-008 wk1=-7.40362e-008 pk1=2.65337e-014 k2=-0.0700206 lk2=3.58404e-008 wk2=1.40211e-008 pk2=-1.41729e-014 k3=0 k3b=0 w0=0 nlx=0 dvt0w=0 dvt1w=0 dvt2w=0 dvt0=0 dvt1=0 
+ dvt2=0 u0=0.0100718 lu0=-1.03686e-009 wu0=-1.00667e-009 pu0=2.36633e-016 ua=1.78672e-009 lua=-5.31135e-016 wua=-4.74914e-016 pua=1.45241e-022 ub=-9.42573e-019 lub=8.36558e-025 wub=2.83937e-025 pub=-1.55429e-031 uc=-2.7142e-010 luc=1.10767e-016 
+ wuc=5.07914e-017 puc=-2.66025e-023 vsat=616436 lvsat=-0.116436 wvsat=0.0399964 pvsat=-3.99964e-008 a0=0.116753 la0=2.64204e-007 wa0=2.49952e-007 pa0=-1.14065e-013 ags=0.0566573 lags=-5.66573e-008 wags=-2.26629e-008 pags=2.26629e-014 b0=0 b1=0 
+ keta=-0.0282549 lketa=2.31327e-009 wketa=1.33697e-008 pketa=-2.27711e-015 a1=0 a2=0.4 rdsw=10 prwg=0.2 prwb=-0.3 wr=1 wint=0 lint=0 dwg=0 dwb=0 voff=-0.211244 lvoff=8.79493e-008 wvoff=1.56624e-008 pvoff=-2.43157e-014 nfactor=11.1853 
+ lnfactor=-4.59264e-006 wnfactor=-3.71033e-006 pnfactor=1.85516e-012 eta0=-0.003669 leta0=2.55311e-009 weta0=1.42773e-009 peta0=-7.55431e-016 etab=0.000711171 letab=-7.11171e-010 wetab=-2.00416e-010 petab=2.00416e-016 pclm=9.207 lpclm=-4.207e-006 
+ wpclm=-1.0278e-006 ppclm=1.0278e-012 pdiblc1=0 pdiblc2=0.194665 lpdiblc2=-9.46653e-008 wpdiblc2=1.59739e-009 ppdiblc2=-1.5974e-015 pdiblcb=0.199414 lpdiblcb=5.85929e-010 wpdiblcb=2.34371e-010 ppdiblcb=-2.34371e-016 drout=0 pscbe1=7.70752e+008 
+ pscbe2=1e-020 pvag=-1 lpvag=1e-006 delta=0.01 ngate=1e+030 dsub=0 cit=-0.0120406 lcit=6.20707e-009 wcit=4.49787e-009 pcit=-2.63289e-015 cdsc=0 cdscd=-0.000152463 lcdscd=1.52463e-010 wcdscd=4.57389e-011 pcdscd=-4.57389e-017 cdscb=0 xpart=0 
+ cgso=2.2653e-010 cgdo=2.2653e-010 cgbo=1e-013 cgsl=0 cgdl=0 ckappa=0.6 cf=0 clc=1e-007 cle=0.6 dlc=0 dwc=0 vfbcv=-0.826159 noff=1 voffcv=0 acde=0.5 moin=15 wln=1 wl=0 wwn=1 ww=0 wwl=0 lln=1 ll=0 lwn=1 lw=0 lwl=0 llc=0 lwc=0 lwlc=0 wlc=0 wwc=0 
+ wwlc=0 alpha0=0 alpha1=0 beta0=30 af=1.1021 kf=1.74179e-023 rsh=3 js=0.0001 jsw=0 cj=0.00150656 mj=0.403022 pb=0.790743 cjsw=1.18641e-010 mjsw=2 tref=27 prt=-149.998 ute=-0.950103 kt1=-0.257006 kt1l=0 kt2=-0.0222175 ua1=1.29549e-010 
+ ub1=-1.58953e-018 uc1=-4.01361e-011 at=-50000 xti=3 tcj=0.00075544 tcjsw=0.0017757 tpb=0.0016635 tpbsw=-0.0013729 elm=5 xl=0 xw=0 ldif=1e-007 hdif=2.7e-007 lmlt=1 wmlt=1 rd=0 rdc=0 rs=0 rsc=0 php=0.8 cjgate=2e-014 n=1 

.model pmos_tkt2.4 pmos level=49 wmax=4e-007 wmin=3e-007 lmax=1e-005 lmin=1e-006 acm=2 version=3.2 mobmod=1 capmod=1 nqsmod=0 binunit=2 binflag=1 tox=5.05e-009 toxm=5.05e-009 xj=1e-007 nch=3.29929e+017 vth0=-0.450058 lvth0=-1.03204e-007 
+ wvth0=2.27213e-008 pvth0=2.76921e-014 vfb=-0.62832 k1=0.408187 lk1=1.59632e-007 wk1=1.94863e-008 pk1=-6.69889e-014 k2=0.0424337 lk2=-7.6614e-008 wk2=-2.7946e-008 pk2=2.77941e-014 k3=0 k3b=0 w0=0 nlx=0 dvt0w=0 dvt1w=0 dvt2w=0 dvt0=0 dvt1=0 dvt2=0 
+ u0=0.00817185 lu0=8.63045e-010 wu0=-1.19623e-011 pu0=-7.58075e-016 ua=4.62042e-010 lua=7.93542e-016 wua=-1.20718e-017 pua=-3.17602e-022 ub=3.24498e-019 lub=-4.30513e-025 wub=-1.485e-025 pub=2.77008e-031 uc=-1.46134e-010 luc=-1.45195e-017 
+ wuc=9.2146e-018 puc=1.49743e-023 vsat=500000 a0=0.990428 la0=-6.09471e-007 wa0=-8.84121e-008 pa0=2.24298e-013 ags=0 b0=0 b1=0 keta=-0.00853487 lketa=-1.74068e-008 wketa=9.98698e-009 pketa=1.10559e-015 a1=0 a2=0.4 rdsw=10 prwg=0.2 prwb=-0.3 wr=1 
+ wint=0 lint=0 dwg=0 dwb=0 voff=-0.0878587 lvoff=-3.54363e-008 wvoff=-2.47595e-008 pvoff=1.61061e-014 nfactor=3.22395 lnfactor=3.36869e-006 wnfactor=-9.11853e-007 pnfactor=-9.43312e-013 eta0=0.00165761 leta0=-2.7735e-009 weta0=-4.60849e-010 
+ peta0=1.13315e-015 etab=0.000829529 letab=-8.29529e-010 wetab=-3.38362e-010 petab=3.38362e-016 pclm=5 pdiblc1=0 pdiblc2=0.1 pdiblcb=0.2 drout=0 pscbe1=7.70752e+008 pscbe2=1e-020 pvag=0 delta=0.01 ngate=1e+030 dsub=0 cit=-0.00606173 
+ lcit=2.28232e-010 wcit=2.62197e-009 pcit=-7.56987e-016 cdsc=0 cdscd=0 cdscb=0 xpart=0 cgso=2.2653e-010 cgdo=2.2653e-010 cgbo=1e-013 cgsl=0 cgdl=0 ckappa=0.6 cf=0 clc=1e-007 cle=0.6 dlc=0 dwc=0 vfbcv=-0.826159 noff=1 voffcv=0 acde=0.5 moin=15 wln=1 
+ wl=0 wwn=1 ww=0 wwl=0 lln=1 ll=0 lwn=1 lw=0 lwl=0 llc=0 lwc=0 lwlc=0 wlc=0 wwc=0 wwlc=0 alpha0=0 alpha1=0 beta0=30 af=1.1021 kf=1.74179e-023 rsh=3 js=0.0001 jsw=0 cj=0.00150656 mj=0.403022 pb=0.790743 cjsw=1.18641e-010 mjsw=2 tref=27 prt=-149.998 
+ ute=-0.950103 kt1=-0.257006 kt1l=0 kt2=-0.0222175 ua1=1.29549e-010 ub1=-1.58953e-018 uc1=-4.01361e-011 at=-50000 xti=3 tcj=0.00075544 tcjsw=0.0017757 tpb=0.0016635 tpbsw=-0.0013729 elm=5 xl=0 xw=0 ldif=1e-007 hdif=2.7e-007 lmlt=1 wmlt=1 rd=0 rdc=0 
+ rs=0 rsc=0 php=0.8 cjgate=2e-014 n=1 

.model pmos_tkt2.5 pmos level=49 wmax=4e-007 wmin=3e-007 lmax=2e-005 lmin=1e-005 acm=2 version=3.2 mobmod=1 capmod=1 nqsmod=0 binunit=2 binflag=1 tox=5.05e-009 toxm=5.05e-009 xj=1e-007 nch=3.29929e+017 vth0=-0.460378 wvth0=2.54905e-008 vfb=-0.62832 
+ k1=0.42415 wk1=1.27875e-008 k2=0.0347723 wk2=-2.51666e-008 k3=0 k3b=0 w0=0 nlx=0 dvt0w=0 dvt1w=0 dvt2w=0 dvt0=0 dvt1=0 dvt2=0 u0=0.00825816 wu0=-8.77698e-011 ua=5.41396e-010 wua=-4.38319e-017 ub=2.81447e-019 wub=-1.208e-025 uc=-1.47586e-010 
+ wuc=1.0712e-017 vsat=500000 a0=0.929481 wa0=-6.59822e-008 ags=0 b0=0 b1=0 keta=-0.0102755 wketa=1.00975e-008 a1=0 a2=0.4 rdsw=10 prwg=0.2 prwb=-0.3 wr=1 wint=0 lint=0 dwg=0 dwb=0 voff=-0.0914024 wvoff=-2.31488e-008 nfactor=3.56082 
+ wnfactor=-1.00618e-006 eta0=0.00138026 weta0=-3.47534e-010 etab=0.000746576 wetab=-3.04526e-010 pclm=5 pdiblc1=0 pdiblc2=0.1 pdiblcb=0.2 drout=0 pscbe1=7.70752e+008 pscbe2=1e-020 pvag=0 delta=0.01 ngate=1e+030 dsub=0 cit=-0.00603891 
+ wcit=2.54627e-009 cdsc=0 cdscd=0 cdscb=0 xpart=0 cgso=2.2653e-010 cgdo=2.2653e-010 cgbo=1e-013 cgsl=0 cgdl=0 ckappa=0.6 cf=0 clc=1e-007 cle=0.6 dlc=0 dwc=0 vfbcv=-0.826159 noff=1 voffcv=0 acde=0.5 moin=15 wln=1 wl=0 wwn=1 ww=0 wwl=0 lln=1 ll=0 
+ lwn=1 lw=0 lwl=0 llc=0 lwc=0 lwlc=0 wlc=0 wwc=0 wwlc=0 alpha0=0 alpha1=0 beta0=30 af=1.1021 kf=1.74179e-023 rsh=3 js=0.0001 jsw=0 cj=0.00150656 mj=0.403022 pb=0.790743 cjsw=1.18641e-010 mjsw=2 tref=27 prt=-149.998 ute=-0.950103 kt1=-0.257006 
+ kt1l=0 kt2=-0.0222175 ua1=1.29549e-010 ub1=-1.58953e-018 uc1=-4.01361e-011 at=-50000 xti=3 tcj=0.00075544 tcjsw=0.0017757 tpb=0.0016635 tpbsw=-0.0013729 elm=5 xl=0 xw=0 ldif=1e-007 hdif=2.7e-007 lmlt=1 wmlt=1 rd=0 rdc=0 rs=0 rsc=0 php=0.8 
+ cjgate=2e-014 n=1 

.model pmos_tkt2.6 pmos level=49 wmax=1e-006 wmin=4e-007 lmax=3e-007 lmin=2.4e-007 acm=2 version=3.2 mobmod=1 capmod=1 nqsmod=0 binunit=2 binflag=1 tox=5.05e-009 toxm=5.05e-009 xj=1e-007 nch=3.29929e+017 vth0=-0.797198 lvth0=6.55164e-008 
+ wvth0=2.60883e-007 pvth0=-5.56501e-014 vfb=-0.62832 k1=0.600533 lk1=-3.23868e-008 wk1=-6.93807e-008 pk1=1.30193e-014 k2=0.0459246 lk2=-2.289e-008 wk2=-1.78192e-008 pk2=4.58824e-015 k3=0 k3b=0 w0=0 nlx=0 dvt0w=0 dvt1w=0 dvt2w=0 dvt0=0 dvt1=0 dvt2=0 
+ u0=0.0134043 lu0=-1.34724e-009 wu0=-5.17036e-009 pu0=1.34059e-015 ua=2.21201e-009 lua=-6.01525e-016 wua=-1.79216e-015 pua=5.41412e-022 ub=1.39135e-018 lub=3.35857e-025 wub=-2.99075e-025 pub=-4.86638e-032 uc=2.65593e-010 luc=-4.05541e-017 
+ wuc=-1.67645e-016 puc=3.62142e-023 vsat=192481 lvsat=0.0116468 wvsat=0.233374 pvsat=-5.40509e-008 a0=-0.519445 la0=3.39993e-008 wa0=8.91523e-007 pa0=-9.08293e-014 ags=0.0201375 lags=-4.12613e-011 wags=-5.50151e-011 pags=1.65045e-017 b0=0 b1=0 
+ keta=0.00760854 lketa=-5.17852e-009 wketa=1.39577e-008 pketa=-1.79487e-015 a1=0 a2=0.4 rdsw=10 prwg=0.2 prwb=-0.3 wr=1 wint=0 lint=0 dwg=0 dwb=0 voff=-0.216448 lvoff=3.80072e-009 wvoff=8.03183e-008 pvoff=-1.20493e-014 nfactor=-4.59351 
+ lnfactor=1.10244e-006 wnfactor=4.59351e-006 pnfactor=-1.10244e-012 eta0=-0.00922745 leta0=3.13393e-009 weta0=2.05579e-009 peta0=-2.70955e-016 etab=-0.00360017 letab=1.65556e-010 wetab=1.03853e-009 petab=-1.34314e-016 pclm=-3.71071 
+ lpclm=1.43128e-006 wpclm=8.18694e-006 ppclm=-1.98331e-012 pdiblc1=0 pdiblc2=0.0121708 lpdiblc2=1.11772e-008 wpdiblc2=-1.16962e-008 ppdiblc2=-2.42133e-015 pdiblcb=-0.738653 lpdiblcb=2.81635e-007 wpdiblcb=1.01507e-006 ppdiblcb=-3.0456e-013 drout=0 
+ pscbe1=7.70752e+008 pscbe2=1e-020 pvag=4.33333 lpvag=-8e-007 wpvag=-3.33333e-006 ppvag=8e-013 delta=0.01 ngate=1e+030 dsub=0 cit=0.00439612 lcit=-8.32408e-010 wcit=-4.51024e-009 pcit=1.12464e-015 cdsc=0 cdscd=-0.000155825 lcdscd=6.28238e-011 
+ wcdscd=9.06468e-011 pcdscd=-2.88316e-017 cdscb=0 xpart=0 cgso=2.2653e-010 cgdo=2.2653e-010 cgbo=1e-013 cgsl=0 cgdl=0 ckappa=0.6 cf=0 clc=1e-007 cle=0.6 dlc=0 dwc=0 vfbcv=-0.826159 noff=1 voffcv=0 acde=0.5 moin=15 wln=1 wl=0 wwn=1 ww=0 wwl=0 lln=1 
+ ll=0 lwn=1 lw=0 lwl=0 llc=0 lwc=0 lwlc=0 wlc=0 wwc=0 wwlc=0 alpha0=0 alpha1=0 beta0=30 af=1.1021 kf=1.74179e-023 rsh=3 js=0.0001 jsw=0 cj=0.00150656 mj=0.403022 pb=0.790743 cjsw=1.18641e-010 mjsw=2 tref=27 prt=-149.998 ute=-0.950103 kt1=-0.257006 
+ kt1l=0 kt2=-0.0222175 ua1=1.29549e-010 ub1=-1.58953e-018 uc1=-4.01361e-011 at=-50000 xti=3 tcj=0.00075544 tcjsw=0.0017757 tpb=0.0016635 tpbsw=-0.0013729 elm=5 xl=0 xw=0 ldif=1e-007 hdif=2.7e-007 lmlt=1 wmlt=1 rd=0 rdc=0 rs=0 rsc=0 php=0.8 
+ cjgate=2e-014 n=1 

.model pmos_tkt2.7 pmos level=49 wmax=1e-006 wmin=4e-007 lmax=5e-007 lmin=3e-007 acm=2 version=3.2 mobmod=1 capmod=1 nqsmod=0 binunit=2 binflag=1 tox=5.05e-009 toxm=5.05e-009 xj=1e-007 nch=3.29929e+017 vth0=-0.46425 lvth0=-3.43679e-008 
+ wvth0=1.58871e-008 pvth0=1.78486e-014 vfb=-0.62832 k1=0.454132 lk1=1.15334e-008 wk1=5.14253e-010 pk1=-7.94924e-015 k2=0.0162829 lk2=-1.39975e-008 wk2=-1.86523e-008 pk2=4.83819e-015 k3=0 k3b=0 w0=0 nlx=0 dvt0w=0 dvt1w=0 dvt2w=0 dvt0=0 dvt1=0 dvt2=0 
+ u0=0.00739897 lu0=4.54367e-010 wu0=-5.90569e-010 pu0=-3.33523e-017 ua=1.42453e-009 lua=-3.65283e-016 wua=-4.49425e-016 pua=1.38592e-022 ub=-5.67769e-019 lub=9.23594e-025 wub=7.57527e-026 pub=-1.61112e-031 uc=-1.30974e-010 luc=7.84162e-017 
+ wuc=-1.13821e-017 puc=-1.06647e-023 vsat=536589 lvsat=-0.0915857 wvsat=-0.149652 pvsat=6.08568e-008 a0=1.13525 la0=-4.6241e-007 wa0=-3.93856e-007 pa0=2.94784e-013 ags=0.0533334 lags=-1e-008 wags=-3.33333e-008 pags=1e-014 b0=0 b1=0 keta=-0.0393505 
+ lketa=8.90919e-009 wketa=7.98019e-009 pketa=-1.61585e-018 a1=0 a2=0.4 rdsw=10 prwg=0.2 prwb=-0.3 wr=1 wint=0 lint=0 dwg=0 dwb=0 voff=-0.0705711 lvoff=-3.99624e-008 wvoff=-2.75036e-008 pvoff=2.02973e-014 nfactor=-1.95528 lnfactor=3.10973e-007 
+ wnfactor=1.95528e-006 pnfactor=-3.10973e-013 eta0=-0.00387747 leta0=1.52894e-009 weta0=3.2008e-010 peta0=2.49758e-016 etab=0.00459168 letab=-2.292e-009 wetab=-1.10403e-009 petab=5.08453e-016 pclm=13.6388 lpclm=-3.77358e-006 wpclm=-5.09302e-006 
+ ppclm=2.00068e-012 pdiblc1=0 pdiblc2=0.0857742 lpdiblc2=-1.09038e-008 wpdiblc2=-3.29745e-008 ppdiblc2=3.96216e-015 pdiblcb=0.199805 lpdiblcb=9.76548e-011 wpdiblcb=1.9531e-010 ppdiblcb=-9.76548e-017 drout=0 pscbe1=7.70752e+008 pscbe2=1e-020 
+ pvag=-4.16667 lpvag=1.75e-006 wpvag=2.66667e-006 ppvag=-1e-012 delta=0.01 ngate=1e+030 dsub=0 cit=0.00462051 lcit=-8.99725e-010 wcit=-3.22512e-009 pcit=7.39107e-016 cdsc=0 cdscd=3.82511e-005 lcdscd=4.60092e-012 wcdscd=-1.14938e-012 
+ pcdscd=-1.29273e-018 cdscb=0 xpart=0 cgso=2.2653e-010 cgdo=2.2653e-010 cgbo=1e-013 cgsl=0 cgdl=0 ckappa=0.6 cf=0 clc=1e-007 cle=0.6 dlc=0 dwc=0 vfbcv=-0.826159 noff=1 voffcv=0 acde=0.5 moin=15 wln=1 wl=0 wwn=1 ww=0 wwl=0 lln=1 ll=0 lwn=1 lw=0 
+ lwl=0 llc=0 lwc=0 lwlc=0 wlc=0 wwc=0 wwlc=0 alpha0=0 alpha1=0 beta0=30 af=1.1021 kf=1.74179e-023 rsh=3 js=0.0001 jsw=0 cj=0.00150656 mj=0.403022 pb=0.790743 cjsw=1.18641e-010 mjsw=2 tref=27 prt=-149.998 ute=-0.950103 kt1=-0.257006 kt1l=0 
+ kt2=-0.0222175 ua1=1.29549e-010 ub1=-1.58953e-018 uc1=-4.01361e-011 at=-50000 xti=3 tcj=0.00075544 tcjsw=0.0017757 tpb=0.0016635 tpbsw=-0.0013729 elm=5 xl=0 xw=0 ldif=1e-007 hdif=2.7e-007 lmlt=1 wmlt=1 rd=0 rdc=0 rs=0 rsc=0 php=0.8 cjgate=2e-014 
+ n=1 

.model pmos_tkt2.8 pmos level=49 wmax=1e-006 wmin=4e-007 lmax=1e-006 lmin=5e-007 acm=2 version=3.2 mobmod=1 capmod=1 nqsmod=0 binunit=2 binflag=1 tox=5.05e-009 toxm=5.05e-009 xj=1e-007 nch=3.29929e+017 vth0=-0.432487 lvth0=-5.02495e-008 
+ wvth0=-7.17779e-009 pvth0=2.93811e-014 vfb=-0.62832 k1=0.432958 lk1=2.21202e-008 wk1=1.05714e-008 pk1=-1.29778e-014 k2=0.0162046 lk2=-1.39583e-008 wk2=-2.0469e-008 pk2=5.74654e-015 k3=0 k3b=0 w0=0 nlx=0 dvt0w=0 dvt1w=0 dvt2w=0 dvt0=0 dvt1=0 dvt2=0 
+ u0=0.0067246 lu0=7.91553e-010 wu0=3.32192e-010 pu0=-4.94733e-016 ua=4.37892e-010 lua=1.28038e-016 wua=6.46163e-017 pua=-1.18428e-022 ub=4.62411e-019 lub=4.08504e-025 wub=-2.78056e-025 pub=1.57922e-032 uc=-1.04346e-010 luc=6.51021e-017 
+ wuc=-1.60383e-017 puc=-8.33665e-024 vsat=646582 lvsat=-0.146582 wvsat=0.0279379 pvsat=-2.79379e-008 a0=0.774176 la0=-2.81872e-007 wa0=-1.30174e-008 pa0=1.04365e-013 ags=0.0333333 wags=-1.33333e-008 b0=0 b1=0 keta=0.0165356 lketa=-1.90339e-008 
+ wketa=-4.54653e-009 pketa=6.26174e-015 a1=0 a2=0.4 rdsw=10 prwg=0.2 prwb=-0.3 wr=1 wint=0 lint=0 dwg=0 dwb=0 voff=-0.170999 lvoff=1.02515e-008 wvoff=-4.35804e-010 pvoff=6.7634e-015 nfactor=-1.27297 lnfactor=-3.01834e-008 wnfactor=1.27297e-006 
+ pnfactor=3.01834e-014 eta0=0.0016719 leta0=-1.24575e-009 weta0=-7.0863e-010 peta0=7.64113e-016 etab=-0.00029384 letab=1.50759e-010 wetab=2.01589e-010 petab=-1.44357e-016 pclm=3.90834 lpclm=1.09166e-006 wpclm=1.09166e-006 ppclm=-1.09166e-012 
+ pdiblc1=0 pdiblc2=0.136033 lpdiblc2=-3.60334e-008 wpdiblc2=2.50502e-008 ppdiblc2=-2.50502e-014 pdiblcb=0.2 drout=0 pscbe1=7.70752e+008 pscbe2=1e-020 pvag=0.666667 lpvag=-6.66667e-007 wpvag=-6.66667e-007 ppvag=6.66667e-013 delta=0.01 ngate=1e+030 
+ dsub=0 cit=0.00133892 lcit=7.41072e-010 wcit=-8.53929e-010 pcit=-4.46488e-016 cdsc=0 cdscd=-4.74529e-005 lcdscd=4.74529e-011 wcdscd=3.73485e-012 pcdscd=-3.73485e-018 cdscb=0 xpart=0 cgso=2.2653e-010 cgdo=2.2653e-010 cgbo=1e-013 cgsl=0 cgdl=0 
+ ckappa=0.6 cf=0 clc=1e-007 cle=0.6 dlc=0 dwc=0 vfbcv=-0.826159 noff=1 voffcv=0 acde=0.5 moin=15 wln=1 wl=0 wwn=1 ww=0 wwl=0 lln=1 ll=0 lwn=1 lw=0 lwl=0 llc=0 lwc=0 lwlc=0 wlc=0 wwc=0 wwlc=0 alpha0=0 alpha1=0 beta0=30 af=1.1021 kf=1.74179e-023 
+ rsh=3 js=0.0001 jsw=0 cj=0.00150656 mj=0.403022 pb=0.790743 cjsw=1.18641e-010 mjsw=2 tref=27 prt=-149.998 ute=-0.950103 kt1=-0.257006 kt1l=0 kt2=-0.0222175 ua1=1.29549e-010 ub1=-1.58953e-018 uc1=-4.01361e-011 at=-50000 xti=3 tcj=0.00075544 
+ tcjsw=0.0017757 tpb=0.0016635 tpbsw=-0.0013729 elm=5 xl=0 xw=0 ldif=1e-007 hdif=2.7e-007 lmlt=1 wmlt=1 rd=0 rdc=0 rs=0 rsc=0 php=0.8 cjgate=2e-014 n=1 

.model pmos_tkt2.9 pmos level=49 wmax=1e-006 wmin=4e-007 lmax=1e-005 lmin=1e-006 acm=2 version=3.2 mobmod=1 capmod=1 nqsmod=0 binunit=2 binflag=1 tox=5.05e-009 toxm=5.05e-009 xj=1e-007 nch=3.29929e+017 vth0=-0.443236 lvth0=-3.95e-008 
+ wvth0=1.99927e-008 pvth0=2.21054e-015 vfb=-0.62832 k1=0.463949 lk1=-8.87057e-009 wk1=-2.81846e-009 pk1=4.12045e-016 k2=0.00508864 lk2=-2.84236e-009 wk2=-1.3008e-008 pk2=-1.71452e-015 k3=0 k3b=0 w0=0 nlx=0 dvt0w=0 dvt1w=0 dvt2w=0 dvt0=0 dvt1=0 
+ dvt2=0 u0=0.00880478 lu0=-1.28863e-009 wu0=-2.65135e-010 pu0=1.02594e-016 ua=7.19856e-010 lua=-1.53926e-016 wua=-1.15197e-016 pua=6.13853e-023 ub=3.9773e-019 lub=4.73185e-025 wub=-1.77793e-025 pub=-8.44708e-032 uc=-9.25745e-011 luc=5.33306e-017 
+ wuc=-1.22092e-017 puc=-1.21657e-023 vsat=500000 a0=0.772007 la0=-2.79703e-007 wa0=-1.04368e-009 pa0=9.23914e-014 ags=0.0333333 wags=-1.33333e-008 b0=0 b1=0 keta=0.0144207 lketa=-1.69189e-008 wketa=8.04768e-010 pketa=9.10447e-016 a1=0 a2=0.4 
+ rdsw=10 prwg=0.2 prwb=-0.213726 lprwb=-8.62745e-008 wprwb=-3.45098e-008 pprwb=3.45098e-014 wr=1 wint=0 lint=0 dwg=0 dwb=0 voff=-0.147295 lvoff=-1.34523e-008 wvoff=-9.84918e-010 pvoff=7.31252e-015 nfactor=-0.629546 lnfactor=-6.73604e-007 
+ wnfactor=6.29546e-007 pnfactor=6.73604e-013 eta0=-0.000144053 leta0=5.70205e-010 weta0=2.59815e-010 peta0=-2.04332e-016 etab=-0.000191765 letab=4.86841e-011 wetab=7.01555e-011 petab=-1.29233e-017 pclm=5 pdiblc1=0 pdiblc2=0.1 pdiblcb=0.2 drout=0 
+ pscbe1=7.70752e+008 pscbe2=1e-020 pvag=0 delta=0.01 ngate=1e+030 dsub=0 cit=0.00170054 lcit=3.79452e-010 wcit=-4.82942e-010 pcit=-8.17475e-016 cdsc=0 cdscd=0 cdscb=0 xpart=0 cgso=2.2653e-010 cgdo=2.2653e-010 cgbo=1e-013 cgsl=0 cgdl=0 ckappa=0.6 
+ cf=0 clc=1e-007 cle=0.6 dlc=0 dwc=0 vfbcv=-0.826159 noff=1 voffcv=0 acde=0.5 moin=15 wln=1 wl=0 wwn=1 ww=0 wwl=0 lln=1 ll=0 lwn=1 lw=0 lwl=0 llc=0 lwc=0 lwlc=0 wlc=0 wwc=0 wwlc=0 alpha0=0 alpha1=0 beta0=30 af=1.1021 kf=1.74179e-023 rsh=3 js=0.0001 
+ jsw=0 cj=0.00150656 mj=0.403022 pb=0.790743 cjsw=1.18641e-010 mjsw=2 tref=27 prt=-149.998 ute=-0.950103 kt1=-0.257006 kt1l=0 kt2=-0.0222175 ua1=1.29549e-010 ub1=-1.58953e-018 uc1=-4.01361e-011 at=-50000 xti=3 tcj=0.00075544 tcjsw=0.0017757 
+ tpb=0.0016635 tpbsw=-0.0013729 elm=5 xl=0 xw=0 ldif=1e-007 hdif=2.7e-007 lmlt=1 wmlt=1 rd=0 rdc=0 rs=0 rsc=0 php=0.8 cjgate=2e-014 n=1 

.model pmos_tkt2.10 pmos level=49 wmax=1e-006 wmin=4e-007 lmax=2e-005 lmin=1e-005 acm=2 version=3.2 mobmod=1 capmod=1 nqsmod=0 binunit=2 binflag=1 tox=5.05e-009 toxm=5.05e-009 xj=1e-007 nch=3.29929e+017 vth0=-0.447186 wvth0=2.02138e-008 vfb=-0.62832 
+ k1=0.463062 wk1=-2.77726e-009 k2=0.0048044 wk2=-1.31794e-008 k3=0 k3b=0 w0=0 nlx=0 dvt0w=0 dvt1w=0 dvt2w=0 dvt0=0 dvt1=0 dvt2=0 u0=0.00867592 wu0=-2.54876e-010 ua=7.04463e-010 wua=-1.09059e-016 ub=4.45048e-019 wub=-1.8624e-025 uc=-8.72414e-011 
+ wuc=-1.34258e-017 vsat=500000 a0=0.744037 wa0=8.19544e-009 ags=0.0333333 wags=-1.33333e-008 b0=0 b1=0 keta=0.0127288 wketa=8.95813e-010 a1=0 a2=0.4 rdsw=10 prwg=0.2 prwb=-0.222353 wprwb=-3.10588e-008 wr=1 wint=0 lint=0 dwg=0 dwb=0 voff=-0.14864 
+ wvoff=-2.53667e-010 nfactor=-0.696906 wnfactor=6.96906e-007 eta0=-8.70325e-005 weta0=2.39382e-010 etab=-0.000186896 wetab=6.88632e-011 pclm=5 pdiblc1=0 pdiblc2=0.1 pdiblcb=0.2 drout=0 pscbe1=7.70752e+008 pscbe2=1e-020 pvag=0 delta=0.01 
+ ngate=1e+030 dsub=0 cit=0.00173848 wcit=-5.6469e-010 cdsc=0 cdscd=0 cdscb=0 xpart=0 cgso=2.2653e-010 cgdo=2.2653e-010 cgbo=1e-013 cgsl=0 cgdl=0 ckappa=0.6 cf=0 clc=1e-007 cle=0.6 dlc=0 dwc=0 vfbcv=-0.826159 noff=1 voffcv=0 acde=0.5 moin=15 wln=1 
+ wl=0 wwn=1 ww=0 wwl=0 lln=1 ll=0 lwn=1 lw=0 lwl=0 llc=0 lwc=0 lwlc=0 wlc=0 wwc=0 wwlc=0 alpha0=0 alpha1=0 beta0=30 af=1.1021 kf=1.74179e-023 rsh=3 js=0.0001 jsw=0 cj=0.00150656 mj=0.403022 pb=0.790743 cjsw=1.18641e-010 mjsw=2 tref=27 prt=-149.998 
+ ute=-0.950103 kt1=-0.257006 kt1l=0 kt2=-0.0222175 ua1=1.29549e-010 ub1=-1.58953e-018 uc1=-4.01361e-011 at=-50000 xti=3 tcj=0.00075544 tcjsw=0.0017757 tpb=0.0016635 tpbsw=-0.0013729 elm=5 xl=0 xw=0 ldif=1e-007 hdif=2.7e-007 lmlt=1 wmlt=1 rd=0 rdc=0 
+ rs=0 rsc=0 php=0.8 cjgate=2e-014 n=1 

.model pmos_tkt2.11 pmos level=49 wmax=1e-005 wmin=1e-006 lmax=3e-007 lmin=2.4e-007 acm=2 version=3.2 mobmod=1 capmod=1 nqsmod=0 binunit=2 binflag=1 tox=5.05e-009 toxm=5.05e-009 xj=1e-007 nch=3.29929e+017 vth0=-0.566142 lvth0=4.16882e-009 
+ wvth0=2.98273e-008 pvth0=5.69745e-015 vfb=-0.62832 k1=0.851692 lk1=-9.0438e-008 wk1=-3.2054e-007 pk1=7.10705e-014 k2=-0.0565962 lk2=2.42953e-009 wk2=8.47016e-008 pk2=-2.07313e-014 k3=0 k3b=0 w0=0 nlx=0 dvt0w=0 dvt1w=0 dvt2w=0 dvt0=0 dvt1=0 dvt2=0 
+ u0=0.00181992 lu0=2.29212e-009 wu0=6.41404e-009 pu0=-2.29877e-015 ua=-2.72237e-009 lua=8.29729e-016 wua=3.14222e-015 pua=-8.89841e-022 ub=9.66913e-019 lub=5.01352e-025 wub=1.25365e-025 pub=-2.14158e-031 uc=-2.79304e-011 luc=5.0877e-017 
+ wuc=1.25879e-016 puc=-5.52169e-023 vsat=406633 lvsat=-0.0326557 wvsat=0.0192221 pvsat=-9.74837e-009 a0=-0.199545 la0=6.37031e-008 wa0=5.71623e-007 pa0=-1.20533e-013 ags=0.0132444 lags=1.62188e-009 wags=6.83808e-009 pags=-1.64664e-015 b0=0 b1=0 
+ keta=-0.0916517 lketa=1.74641e-008 wketa=1.13218e-007 pketa=-2.44375e-014 a1=0 a2=0.4 rdsw=10 prwg=0.2 prwb=-0.3 wr=1 wint=0 lint=0 dwg=0 dwb=0 voff=-0.0817371 lvoff=-9.08856e-009 wvoff=-5.43927e-008 pvoff=8.39998e-016 nfactor=-0.801161 
+ lnfactor=2.40348e-007 wnfactor=8.01161e-007 pnfactor=-2.40348e-013 eta0=-0.0249601 leta0=8.23484e-009 weta0=1.77884e-008 peta0=-5.37187e-015 etab=0.00239398 letab=-1.16607e-009 wetab=-4.95563e-009 petab=1.19732e-015 pclm=4.37664 
+ lpclm=-7.93474e-007 wpclm=9.96018e-008 ppclm=2.41442e-013 pdiblc1=0 pdiblc2=0.14384 lpdiblc2=-3.38073e-008 wpdiblc2=-1.43365e-007 ppdiblc2=4.25631e-014 pdiblcb=0.191509 lpdiblcb=2.54723e-009 wpdiblcb=8.49075e-008 ppdiblcb=-2.54723e-014 drout=0 
+ pscbe1=7.70752e+008 pscbe2=1e-020 pvag=1 delta=0.01 ngate=1e+030 dsub=0 cit=0.00172914 lcit=-3.04451e-011 wcit=-1.84325e-009 pcit=3.2268e-016 cdsc=0 cdscd=0.000199697 lcdscd=-4.92933e-011 wcdscd=-2.64876e-010 pcdscd=8.32855e-017 cdscb=0 xpart=0 
+ cgso=2.2653e-010 cgdo=2.2653e-010 cgbo=1e-013 cgsl=0 cgdl=0 ckappa=0.6 cf=0 clc=1e-007 cle=0.6 dlc=0 dwc=0 vfbcv=-0.826159 noff=1 voffcv=0 acde=0.5 moin=15 wln=1 wl=0 wwn=1 ww=0 wwl=0 lln=1 ll=0 lwn=1 lw=0 lwl=0 llc=0 lwc=0 lwlc=0 wlc=0 wwc=0 
+ wwlc=0 alpha0=0 alpha1=0 beta0=30 af=1.1021 kf=1.74179e-023 rsh=3 js=0.0001 jsw=0 cj=0.00150656 mj=0.403022 pb=0.790743 cjsw=1.18641e-010 mjsw=2 tref=27 prt=-149.998 ute=-0.950103 kt1=-0.257006 kt1l=0 kt2=-0.0222175 ua1=1.29549e-010 
+ ub1=-1.58953e-018 uc1=-4.01361e-011 at=-50000 xti=3 tcj=0.00075544 tcjsw=0.0017757 tpb=0.0016635 tpbsw=-0.0013729 elm=5 xl=0 xw=0 ldif=1e-007 hdif=2.7e-007 lmlt=1 wmlt=1 rd=0 rdc=0 rs=0 rsc=0 php=0.8 cjgate=2e-014 n=1 

.model pmos_tkt2.12 pmos level=49 wmax=1e-005 wmin=1e-006 lmax=5e-007 lmin=3e-007 acm=2 version=3.2 mobmod=1 capmod=1 nqsmod=0 binunit=2 binflag=1 tox=5.05e-009 toxm=5.05e-009 xj=1e-007 nch=3.29929e+017 vth0=-0.45473 lvth0=-2.9255e-008 
+ wvth0=6.36662e-009 pvth0=1.27356e-014 vfb=-0.62832 k1=0.426955 lk1=3.69833e-008 wk1=2.76918e-008 pk1=-3.33992e-014 k2=0.0334634 lk2=-2.45884e-008 wk2=-3.58329e-008 pk2=1.54291e-014 k3=0 k3b=0 w0=0 nlx=0 dvt0w=0 dvt1w=0 dvt2w=0 dvt0=0 dvt1=0 dvt2=0 
+ u0=0.00766224 lu0=5.39424e-010 wu0=-8.5384e-010 pu0=-1.18409e-016 ua=1.0951e-009 lua=-3.15513e-016 wua=-1.19987e-016 pua=8.88215e-023 ub=-7.01331e-021 lub=7.9353e-025 wub=-4.85003e-025 pub=-3.10477e-032 uc=-8.8667e-011 luc=6.9098e-017 
+ wuc=-5.36894e-017 puc=-1.34643e-024 vsat=851807 lvsat=-0.166208 wvsat=-0.464869 pvsat=1.35479e-007 a0=0.671883 la0=-1.97726e-007 wa0=6.95118e-008 pa0=3.01003e-014 ags=0.0220239 lags=-1.01196e-009 wags=-2.02392e-009 pags=1.01196e-015 b0=0 b1=0 
+ keta=-0.00772459 lketa=-7.71403e-009 wketa=-2.36457e-008 pketa=1.66216e-014 a1=0 a2=0.4 rdsw=10 prwg=0.2 prwb=-0.3 wr=1 wint=0 lint=0 dwg=0 dwb=0 voff=-0.155678 lvoff=1.30938e-008 wvoff=5.76034e-008 pvoff=-3.27588e-014 nfactor=0 eta0=-0.00338606 
+ leta0=1.76263e-009 weta0=-1.71329e-010 peta0=1.6061e-017 etab=0.000536796 letab=-6.08918e-010 wetab=2.95085e-009 petab=-1.17463e-015 pclm=9.90242 lpclm=-2.45121e-006 wpclm=-1.35661e-006 ppclm=6.78307e-013 pdiblc1=0 pdiblc2=0.220244 
+ lpdiblc2=-5.67286e-008 wpdiblc2=-1.67445e-007 ppdiblc2=4.9787e-014 pdiblcb=0.2 drout=0 pscbe1=7.70752e+008 pscbe2=1e-020 pvag=-1.5 lpvag=7.5e-007 delta=0.01 ngate=1e+030 dsub=0 cit=0.000819814 lcit=2.42352e-010 wcit=5.75578e-010 pcit=-4.02969e-016 
+ cdsc=0 cdscd=-2.59025e-005 lcdscd=1.83866e-011 wcdscd=6.30042e-011 pcdscd=-1.50784e-017 cdscb=0 xpart=0 cgso=2.2653e-010 cgdo=2.2653e-010 cgbo=1e-013 cgsl=0 cgdl=0 ckappa=0.6 cf=0 clc=1e-007 cle=0.6 dlc=0 dwc=0 vfbcv=-0.826159 noff=1 voffcv=0 
+ acde=0.5 moin=15 wln=1 wl=0 wwn=1 ww=0 wwl=0 lln=1 ll=0 lwn=1 lw=0 lwl=0 llc=0 lwc=0 lwlc=0 wlc=0 wwc=0 wwlc=0 alpha0=0 alpha1=0 beta0=30 af=1.1021 kf=1.74179e-023 rsh=3 js=0.0001 jsw=0 cj=0.00150656 mj=0.403022 pb=0.790743 cjsw=1.18641e-010 
+ mjsw=2 tref=27 prt=-149.998 ute=-0.950103 kt1=-0.257006 kt1l=0 kt2=-0.0222175 ua1=1.29549e-010 ub1=-1.58953e-018 uc1=-4.01361e-011 at=-50000 xti=3 tcj=0.00075544 tcjsw=0.0017757 tpb=0.0016635 tpbsw=-0.0013729 elm=5 xl=0 xw=0 ldif=1e-007 
+ hdif=2.7e-007 lmlt=1 wmlt=1 rd=0 rdc=0 rs=0 rsc=0 php=0.8 cjgate=2e-014 n=1 

.model pmos_tkt2.13 pmos level=49 wmax=1e-005 wmin=1e-006 lmax=1e-006 lmin=5e-007 acm=2 version=3.2 mobmod=1 capmod=1 nqsmod=0 binunit=2 binflag=1 tox=5.05e-009 toxm=5.05e-009 xj=1e-007 nch=3.29929e+017 vth0=-0.458425 lvth0=-2.74074e-008 
+ wvth0=1.87599e-008 pvth0=6.53903e-015 vfb=-0.62832 k1=0.486548 lk1=7.18684e-009 wk1=-4.30177e-008 pk1=1.95556e-015 k2=-0.0047544 lk2=-5.47945e-009 wk2=4.90005e-010 pk2=-2.73236e-015 k3=0 k3b=0 w0=0 nlx=0 dvt0w=0 dvt1w=0 dvt2w=0 dvt0=0 dvt1=0 
+ dvt2=0 u0=0.00862235 lu0=5.93721e-011 wu0=-1.56556e-009 pu0=2.37448e-016 ua=8.85709e-010 lua=-2.10819e-016 wua=-3.83201e-016 pua=2.20428e-022 ub=3.41507e-019 lub=6.19269e-025 wub=-1.57152e-025 pub=-1.94973e-031 uc=-1.05014e-010 luc=7.72716e-017 
+ wuc=-1.53701e-017 puc=-2.05061e-023 vsat=480609 lvsat=0.0193911 wvsat=0.193911 pvsat=-1.93911e-007 a0=0.680921 la0=-2.02245e-007 wa0=8.02371e-008 pa0=2.47377e-014 ags=0.02 b0=0 b1=0 keta=0.00981639 lketa=-1.64845e-008 wketa=2.17267e-009 
+ pketa=3.7124e-015 a1=0 a2=0.4 rdsw=10 prwg=0.2 prwb=-0.3 wr=1 wint=0 lint=0 dwg=0 dwb=0 voff=-0.100121 lvoff=-1.46847e-008 wvoff=-7.13133e-008 pvoff=3.16995e-014 nfactor=0.335326 lnfactor=-1.67663e-007 wnfactor=-3.35326e-007 pnfactor=1.67663e-013 
+ eta0=0.000642356 leta0=-2.51574e-010 weta0=3.20915e-010 peta0=-2.30061e-016 etab=0.000533291 letab=-6.07165e-010 wetab=-6.25542e-010 petab=6.13567e-016 pclm=5 pdiblc1=0 pdiblc2=0.0932129 lpdiblc2=6.78706e-009 wpdiblc2=6.78706e-008 
+ ppdiblc2=-6.78706e-014 pdiblcb=0.2 drout=0 pscbe1=7.70752e+008 pscbe2=1e-020 pvag=0 delta=0.01 ngate=1e+030 dsub=0 cit=0.00137234 lcit=-3.39103e-011 wcit=-8.87349e-010 pcit=3.28494e-016 cdsc=0 cdscd=1.50168e-005 lcdscd=-2.07308e-012 
+ wcdscd=-5.87349e-011 pcdscd=4.57911e-017 cdscb=0 xpart=0 cgso=2.2653e-010 cgdo=2.2653e-010 cgbo=1e-013 cgsl=0 cgdl=0 ckappa=0.6 cf=0 clc=1e-007 cle=0.6 dlc=0 dwc=0 vfbcv=-0.826159 noff=1 voffcv=0 acde=0.5 moin=15 wln=1 wl=0 wwn=1 ww=0 wwl=0 lln=1 
+ ll=0 lwn=1 lw=0 lwl=0 llc=0 lwc=0 lwlc=0 wlc=0 wwc=0 wwlc=0 alpha0=0 alpha1=0 beta0=30 af=1.1021 kf=1.74179e-023 rsh=3 js=0.0001 jsw=0 cj=0.00150656 mj=0.403022 pb=0.790743 cjsw=1.18641e-010 mjsw=2 tref=27 prt=-149.998 ute=-0.950103 kt1=-0.257006 
+ kt1l=0 kt2=-0.0222175 ua1=1.29549e-010 ub1=-1.58953e-018 uc1=-4.01361e-011 at=-50000 xti=3 tcj=0.00075544 tcjsw=0.0017757 tpb=0.0016635 tpbsw=-0.0013729 elm=5 xl=0 xw=0 ldif=1e-007 hdif=2.7e-007 lmlt=1 wmlt=1 rd=0 rdc=0 rs=0 rsc=0 php=0.8 
+ cjgate=2e-014 n=1 

.model pmos_tkt2.14 pmos level=49 wmax=1e-005 wmin=1e-006 lmax=1e-005 lmin=1e-006 acm=2 version=3.2 mobmod=1 capmod=1 nqsmod=0 binunit=2 binflag=1 tox=5.05e-009 toxm=5.05e-009 xj=1e-007 nch=3.29929e+017 vth0=-0.43417 lvth0=-5.16625e-008 
+ wvth0=1.09258e-008 pvth0=1.43731e-014 vfb=-0.62832 k1=0.508258 lk1=-1.45239e-008 wk1=-4.71274e-008 pk1=6.06532e-015 k2=-0.00901429 lk2=-1.21956e-009 wk2=1.09497e-009 pk2=-3.33732e-015 k3=0 k3b=0 w0=0 nlx=0 dvt0w=0 dvt1w=0 dvt2w=0 dvt0=0 dvt1=0 
+ dvt2=0 u0=0.00949313 lu0=-8.11411e-010 wu0=-9.53484e-010 pu0=-3.74623e-016 ua=6.42503e-010 lua=3.23869e-017 wua=-3.78446e-017 pua=-1.24928e-022 ub=5.68239e-019 lub=3.92537e-025 wub=-3.48302e-025 pub=-3.82284e-033 uc=-7.96577e-011 luc=5.19151e-017 
+ wuc=-2.5126e-017 puc=-1.07502e-023 vsat=500000 a0=0.681057 la0=-2.0238e-007 wa0=8.99064e-008 pa0=1.50684e-014 ags=0.02 b0=0 b1=0 keta=0.0120469 lketa=-1.87151e-008 wketa=3.17849e-009 pketa=2.70658e-015 a1=0 a2=0.4 rdsw=10 prwg=0.2 prwb=-0.155536 
+ lprwb=-1.44464e-007 wprwb=-9.2699e-008 pprwb=9.2699e-014 wr=1 wint=0 lint=0 dwg=0 dwb=0 voff=-0.116757 lvoff=1.95133e-009 wvoff=-3.15227e-008 pvoff=-8.0911e-015 nfactor=0.0379668 lnfactor=1.29696e-007 wnfactor=-3.79668e-008 pnfactor=-1.29696e-013 
+ eta0=-6.22288e-005 leta0=4.53011e-010 weta0=1.77991e-010 peta0=-8.7137e-017 etab=-0.000125695 letab=5.18204e-011 wetab=4.08553e-012 petab=-1.60596e-017 pclm=5 pdiblc1=0 pdiblc2=0.1 pdiblcb=0.2 drout=0 pscbe1=7.70752e+008 pscbe2=1e-020 pvag=0 
+ delta=0.01 ngate=1e+030 dsub=0 cit=0.00112335 lcit=2.15076e-010 wcit=9.42437e-011 pcit=-6.53099e-016 cdsc=0 cdscd=2.31917e-005 lcdscd=-1.02479e-011 wcdscd=-2.31917e-011 pcdscd=1.02479e-017 cdscb=0 xpart=0 cgso=2.2653e-010 cgdo=2.2653e-010 
+ cgbo=1e-013 cgsl=0 cgdl=0 ckappa=0.6 cf=0 clc=1e-007 cle=0.6 dlc=0 dwc=0 vfbcv=-0.826159 noff=1 voffcv=0 acde=0.5 moin=15 wln=1 wl=0 wwn=1 ww=0 wwl=0 lln=1 ll=0 lwn=1 lw=0 lwl=0 llc=0 lwc=0 lwlc=0 wlc=0 wwc=0 wwlc=0 alpha0=0 alpha1=0 beta0=30 
+ af=1.1021 kf=1.74179e-023 rsh=3 js=0.0001 jsw=0 cj=0.00150656 mj=0.403022 pb=0.790743 cjsw=1.18641e-010 mjsw=2 tref=27 prt=-149.998 ute=-0.950103 kt1=-0.257006 kt1l=0 kt2=-0.0222175 ua1=1.29549e-010 ub1=-1.58953e-018 uc1=-4.01361e-011 at=-50000 
+ xti=3 tcj=0.00075544 tcjsw=0.0017757 tpb=0.0016635 tpbsw=-0.0013729 elm=5 xl=0 xw=0 ldif=1e-007 hdif=2.7e-007 lmlt=1 wmlt=1 rd=0 rdc=0 rs=0 rsc=0 php=0.8 cjgate=2e-014 n=1 

.model pmos_tkt2.15 pmos level=49 wmax=1e-005 wmin=1e-006 lmax=2e-005 lmin=1e-005 acm=2 version=3.2 mobmod=1 capmod=1 nqsmod=0 binunit=2 binflag=1 tox=5.05e-009 toxm=5.05e-009 xj=1e-007 nch=3.29929e+017 vth0=-0.439336 wvth0=1.23631e-008 vfb=-0.62832 
+ k1=0.506806 wk1=-4.65209e-008 k2=-0.00913624 wk2=7.61234e-010 k3=0 k3b=0 w0=0 nlx=0 dvt0w=0 dvt1w=0 dvt2w=0 dvt0=0 dvt1=0 dvt2=0 u0=0.00941199 wu0=-9.90947e-010 ua=6.45742e-010 wua=-5.03373e-017 ub=6.07493e-019 wub=-3.48685e-025 uc=-7.44662e-011 
+ wuc=-2.6201e-017 vsat=500000 a0=0.660819 wa0=9.14133e-008 ags=0.02 b0=0 b1=0 keta=0.0101754 wketa=3.44914e-009 a1=0 a2=0.4 rdsw=10 prwg=0.2 prwb=-0.169983 wprwb=-8.34291e-008 wr=1 wint=0 lint=0 dwg=0 dwb=0 voff=-0.116562 wvoff=-3.23318e-008 
+ nfactor=0.0509365 wnfactor=-5.09364e-008 eta0=-1.69277e-005 weta0=1.69277e-010 etab=-0.000120513 wetab=2.47957e-012 pclm=5 pdiblc1=0 pdiblc2=0.1 pdiblcb=0.2 drout=0 pscbe1=7.70752e+008 pscbe2=1e-020 pvag=0 delta=0.01 ngate=1e+030 dsub=0 
+ cit=0.00114486 wcit=2.89339e-011 cdsc=0 cdscd=2.21669e-005 wcdscd=-2.21669e-011 cdscb=0 xpart=0 cgso=2.2653e-010 cgdo=2.2653e-010 cgbo=1e-013 cgsl=0 cgdl=0 ckappa=0.6 cf=0 clc=1e-007 cle=0.6 dlc=0 dwc=0 vfbcv=-0.826159 noff=1 voffcv=0 acde=0.5 
+ moin=15 wln=1 wl=0 wwn=1 ww=0 wwl=0 lln=1 ll=0 lwn=1 lw=0 lwl=0 llc=0 lwc=0 lwlc=0 wlc=0 wwc=0 wwlc=0 alpha0=0 alpha1=0 beta0=30 af=1.1021 kf=1.74179e-023 rsh=3 js=0.0001 jsw=0 cj=0.00150656 mj=0.403022 pb=0.790743 cjsw=1.18641e-010 mjsw=2 tref=27 
+ prt=-149.998 ute=-0.950103 kt1=-0.257006 kt1l=0 kt2=-0.0222175 ua1=1.29549e-010 ub1=-1.58953e-018 uc1=-4.01361e-011 at=-50000 xti=3 tcj=0.00075544 tcjsw=0.0017757 tpb=0.0016635 tpbsw=-0.0013729 elm=5 xl=0 xw=0 ldif=1e-007 hdif=2.7e-007 lmlt=1 
+ wmlt=1 rd=0 rdc=0 rs=0 rsc=0 php=0.8 cjgate=2e-014 n=1 

.model pmos_tkt2.16 pmos level=49 wmax=0.0001 wmin=1e-005 lmax=3e-007 lmin=2.4e-007 acm=2 version=3.2 mobmod=1 capmod=1 nqsmod=0 binunit=2 binflag=1 tox=5.05e-009 toxm=5.05e-009 xj=1e-007 nch=3.29929e+017 vth0=-0.56316 lvth0=4.73857e-009 
+ vfb=-0.62832 k1=0.819638 lk1=-8.3331e-008 k2=-0.048126 lk2=3.56398e-010 k3=0 k3b=0 w0=0 nlx=0 dvt0w=0 dvt1w=0 dvt2w=0 dvt0=0 dvt1=0 dvt2=0 u0=0.00246132 lu0=2.06225e-009 ua=-2.40815e-009 lua=7.40744e-016 ub=9.7945e-019 lub=4.79936e-025 
+ uc=-1.53425e-011 luc=4.53553e-017 vsat=408555 lvsat=-0.0336306 a0=-0.142383 la0=5.16497e-008 ags=0.0139283 lags=1.45722e-009 b0=0 b1=0 keta=-0.0803299 lketa=1.50204e-008 a1=0 a2=0.4 rdsw=10 prwg=0.2 prwb=-0.3 wr=1 wint=0 lint=0 dwg=0 dwb=0 
+ voff=-0.0871764 lvoff=-9.00456e-009 nfactor=-0.721044 lnfactor=2.16313e-007 eta0=-0.0231812 leta0=7.69765e-009 etab=0.00189842 letab=-1.04634e-009 pclm=4.38659 lpclm=-7.6933e-007 pdiblc1=0 pdiblc2=0.129503 lpdiblc2=-2.95509e-008 pdiblcb=0.2 
+ drout=0 pscbe1=7.70752e+008 pscbe2=1e-020 pvag=1 delta=0.01 ngate=1e+030 dsub=0 cit=0.00154481 lcit=1.82292e-012 cdsc=0 cdscd=0.00017321 lcdscd=-4.09648e-011 cdscb=0 xpart=0 cgso=2.2653e-010 cgdo=2.2653e-010 cgbo=1e-013 cgsl=0 cgdl=0 ckappa=0.6 
+ cf=0 clc=1e-007 cle=0.6 dlc=0 dwc=0 vfbcv=-0.826159 noff=1 voffcv=0 acde=0.5 moin=15 wln=1 wl=0 wwn=1 ww=0 wwl=0 lln=1 ll=0 lwn=1 lw=0 lwl=0 llc=0 lwc=0 lwlc=0 wlc=0 wwc=0 wwlc=0 alpha0=0 alpha1=0 beta0=30 af=1.1021 kf=1.74179e-023 rsh=3 js=0.0001 
+ jsw=0 cj=0.00150656 mj=0.403022 pb=0.790743 cjsw=1.18641e-010 mjsw=2 tref=27 prt=-149.998 ute=-0.950103 kt1=-0.257006 kt1l=0 kt2=-0.0222175 ua1=1.29549e-010 ub1=-1.58953e-018 uc1=-4.01361e-011 at=-50000 xti=3 tcj=0.00075544 tcjsw=0.0017757 
+ tpb=0.0016635 tpbsw=-0.0013729 elm=5 xl=0 xw=0 ldif=1e-007 hdif=2.7e-007 lmlt=1 wmlt=1 rd=0 rdc=0 rs=0 rsc=0 php=0.8 cjgate=2e-014 n=1 

.model pmos_tkt2.17 pmos level=49 wmax=0.0001 wmin=1e-005 lmax=5e-007 lmin=3e-007 acm=2 version=3.2 mobmod=1 capmod=1 nqsmod=0 binunit=2 binflag=1 tox=5.05e-009 toxm=5.05e-009 xj=1e-007 nch=3.29929e+017 vth0=-0.454093 lvth0=-2.79814e-008 
+ vfb=-0.62832 k1=0.429724 lk1=3.36434e-008 k2=0.0298801 lk2=-2.30455e-008 k3=0 k3b=0 w0=0 nlx=0 dvt0w=0 dvt1w=0 dvt2w=0 dvt0=0 dvt1=0 dvt2=0 u0=0.00757686 lu0=5.27584e-010 ua=1.0831e-009 lua=-3.06631e-016 ub=-5.55135e-020 lub=7.90425e-025 
+ uc=-9.40359e-011 luc=6.89633e-017 vsat=805320 lvsat=-0.15266 a0=0.678834 la0=-1.94716e-007 ags=0.0218215 lags=-9.10762e-010 b0=0 b1=0 keta=-0.0100892 lketa=-6.05187e-009 a1=0 a2=0.4 rdsw=10 prwg=0.2 prwb=-0.3 wr=1 wint=0 lint=0 dwg=0 dwb=0 
+ voff=-0.149918 lvoff=9.81788e-009 nfactor=0 eta0=-0.00340319 leta0=1.76424e-009 etab=0.000831881 letab=-7.2638e-010 pclm=9.76676 lpclm=-2.38338e-006 pdiblc1=0 pdiblc2=0.2035 lpdiblc2=-5.17499e-008 pdiblcb=0.2 drout=0 pscbe1=7.70752e+008 
+ pscbe2=1e-020 pvag=-1.5 lpvag=7.5e-007 delta=0.01 ngate=1e+030 dsub=0 cit=0.000877372 lcit=2.02055e-010 cdsc=0 cdscd=-1.96021e-005 lcdscd=1.68788e-011 cdscb=0 xpart=0 cgso=2.2653e-010 cgdo=2.2653e-010 cgbo=1e-013 cgsl=0 cgdl=0 ckappa=0.6 cf=0 
+ clc=1e-007 cle=0.6 dlc=0 dwc=0 vfbcv=-0.826159 noff=1 voffcv=0 acde=0.5 moin=15 wln=1 wl=0 wwn=1 ww=0 wwl=0 lln=1 ll=0 lwn=1 lw=0 lwl=0 llc=0 lwc=0 lwlc=0 wlc=0 wwc=0 wwlc=0 alpha0=0 alpha1=0 beta0=30 af=1.1021 kf=1.74179e-023 rsh=3 js=0.0001 
+ jsw=0 cj=0.00150656 mj=0.403022 pb=0.790743 cjsw=1.18641e-010 mjsw=2 tref=27 prt=-149.998 ute=-0.950103 kt1=-0.257006 kt1l=0 kt2=-0.0222175 ua1=1.29549e-010 ub1=-1.58953e-018 uc1=-4.01361e-011 at=-50000 xti=3 tcj=0.00075544 tcjsw=0.0017757 
+ tpb=0.0016635 tpbsw=-0.0013729 elm=5 xl=0 xw=0 ldif=1e-007 hdif=2.7e-007 lmlt=1 wmlt=1 rd=0 rdc=0 rs=0 rsc=0 php=0.8 cjgate=2e-014 n=1 

.model pmos_tkt2.18 pmos level=49 wmax=0.0001 wmin=1e-005 lmax=1e-006 lmin=5e-007 acm=2 version=3.2 mobmod=1 capmod=1 nqsmod=0 binunit=2 binflag=1 tox=5.05e-009 toxm=5.05e-009 xj=1e-007 nch=3.29929e+017 vth0=-0.456549 lvth0=-2.67535e-008 
+ vfb=-0.62832 k1=0.482246 lk1=7.38239e-009 k2=-0.0047054 lk2=-5.75268e-009 k3=0 k3b=0 w0=0 nlx=0 dvt0w=0 dvt1w=0 dvt2w=0 dvt0=0 dvt1=0 dvt2=0 u0=0.00846579 lu0=8.31169e-011 ua=8.47389e-010 lua=-1.88776e-016 ub=3.25792e-019 lub=5.99772e-025 
+ uc=-1.06551e-010 luc=7.52209e-017 vsat=500000 a0=0.688945 la0=-1.99771e-007 ags=0.02 b0=0 b1=0 keta=0.0100337 lketa=-1.61133e-008 a1=0 a2=0.4 rdsw=10 prwg=0.2 prwb=-0.3 wr=1 wint=0 lint=0 dwg=0 dwb=0 voff=-0.107253 lvoff=-1.15147e-008 
+ nfactor=0.301793 lnfactor=-1.50897e-007 eta0=0.000674448 leta0=-2.7458e-010 etab=0.000470737 letab=-5.45808e-010 pclm=5 pdiblc1=0 pdiblc2=0.1 pdiblcb=0.2 drout=0 pscbe1=7.70752e+008 pscbe2=1e-020 pvag=0 delta=0.01 ngate=1e+030 dsub=0 cit=0.0012836 
+ lcit=-1.06089e-012 cdsc=0 cdscd=9.14335e-006 lcdscd=2.50603e-012 cdscb=0 xpart=0 cgso=2.2653e-010 cgdo=2.2653e-010 cgbo=1e-013 cgsl=0 cgdl=0 ckappa=0.6 cf=0 clc=1e-007 cle=0.6 dlc=0 dwc=0 vfbcv=-0.826159 noff=1 voffcv=0 acde=0.5 moin=15 wln=1 wl=0 
+ wwn=1 ww=0 wwl=0 lln=1 ll=0 lwn=1 lw=0 lwl=0 llc=0 lwc=0 lwlc=0 wlc=0 wwc=0 wwlc=0 alpha0=0 alpha1=0 beta0=30 af=1.1021 kf=1.74179e-023 rsh=3 js=0.0001 jsw=0 cj=0.00150656 mj=0.403022 pb=0.790743 cjsw=1.18641e-010 mjsw=2 tref=27 prt=-149.998 
+ ute=-0.950103 kt1=-0.257006 kt1l=0 kt2=-0.0222175 ua1=1.29549e-010 ub1=-1.58953e-018 uc1=-4.01361e-011 at=-50000 xti=3 tcj=0.00075544 tcjsw=0.0017757 tpb=0.0016635 tpbsw=-0.0013729 elm=5 xl=0 xw=0 ldif=1e-007 hdif=2.7e-007 lmlt=1 wmlt=1 rd=0 rdc=0 
+ rs=0 rsc=0 php=0.8 cjgate=2e-014 n=1 

.model pmos_tkt2.19 pmos level=49 wmax=0.0001 wmin=1e-005 lmax=1e-005 lmin=1e-006 acm=2 version=3.2 mobmod=1 capmod=1 nqsmod=0 binunit=2 binflag=1 tox=5.05e-009 toxm=5.05e-009 xj=1e-007 nch=3.29929e+017 vth0=-0.433077 lvth0=-5.02252e-008 
+ vfb=-0.62832 k1=0.503545 lk1=-1.39173e-008 k2=-0.00890479 lk2=-1.55329e-009 k3=0 k3b=0 w0=0 nlx=0 dvt0w=0 dvt1w=0 dvt2w=0 dvt0=0 dvt1=0 dvt2=0 u0=0.00939778 lu0=-8.48874e-010 ua=6.38719e-010 lua=1.98941e-017 ub=5.33409e-019 lub=3.92155e-025 
+ uc=-8.21703e-011 luc=5.084e-017 vsat=500000 a0=0.690047 la0=-2.00873e-007 ags=0.02 b0=0 b1=0 keta=0.0123648 lketa=-1.84444e-008 a1=0 a2=0.4 rdsw=10 prwg=0.2 prwb=-0.164806 lprwb=-1.35194e-007 wr=1 wint=0 lint=0 dwg=0 dwb=0 voff=-0.11991 
+ lvoff=1.14222e-009 nfactor=0.0341702 lnfactor=1.16726e-007 eta0=-4.44297e-005 leta0=4.44297e-010 etab=-0.000125286 letab=5.02144e-011 pclm=5 pdiblc1=0 pdiblc2=0.1 pdiblcb=0.2 drout=0 pscbe1=7.70752e+008 pscbe2=1e-020 pvag=0 delta=0.01 ngate=1e+030 
+ dsub=0 cit=0.00113278 lcit=1.49766e-010 cdsc=0 cdscd=2.08725e-005 lcdscd=-9.22312e-012 cdscb=0 xpart=0 cgso=2.2653e-010 cgdo=2.2653e-010 cgbo=1e-013 cgsl=0 cgdl=0 ckappa=0.6 cf=0 clc=1e-007 cle=0.6 dlc=0 dwc=0 vfbcv=-0.826159 noff=1 voffcv=0 
+ acde=0.5 moin=15 wln=1 wl=0 wwn=1 ww=0 wwl=0 lln=1 ll=0 lwn=1 lw=0 lwl=0 llc=0 lwc=0 lwlc=0 wlc=0 wwc=0 wwlc=0 alpha0=0 alpha1=0 beta0=30 af=1.1021 kf=1.74179e-023 rsh=3 js=0.0001 jsw=0 cj=0.00150656 mj=0.403022 pb=0.790743 cjsw=1.18641e-010 
+ mjsw=2 tref=27 prt=-149.998 ute=-0.950103 kt1=-0.257006 kt1l=0 kt2=-0.0222175 ua1=1.29549e-010 ub1=-1.58953e-018 uc1=-4.01361e-011 at=-50000 xti=3 tcj=0.00075544 tcjsw=0.0017757 tpb=0.0016635 tpbsw=-0.0013729 elm=5 xl=0 xw=0 ldif=1e-007 
+ hdif=2.7e-007 lmlt=1 wmlt=1 rd=0 rdc=0 rs=0 rsc=0 php=0.8 cjgate=2e-014 n=1 

.model pmos_tkt2.20 pmos level=49 wmax=0.0001 wmin=1e-005 lmax=2e-005 lmin=1e-005 acm=2 version=3.2 mobmod=1 capmod=1 nqsmod=0 binunit=2 binflag=1 tox=5.05e-009 toxm=5.05e-009 xj=1e-007 nch=3.29929e+017 vth0=-0.438099 vfb=-0.62832 k1=0.502154 
+ k2=-0.00906012 k3=0 k3b=0 w0=0 nlx=0 dvt0w=0 dvt1w=0 dvt2w=0 dvt0=0 dvt1=0 dvt2=0 u0=0.0093129 ua=6.40708e-010 ub=5.72625e-019 uc=-7.70863e-011 vsat=500000 a0=0.66996 ags=0.02 b0=0 b1=0 keta=0.0105204 a1=0 a2=0.4 rdsw=10 prwg=0.2 prwb=-0.178326 
+ wr=1 wint=0 lint=0 dwg=0 dwb=0 voff=-0.119795 nfactor=0.0458428 eta0=0 etab=-0.000120265 pclm=5 pdiblc1=0 pdiblc2=0.1 pdiblcb=0.2 drout=0 pscbe1=7.70752e+008 pscbe2=1e-020 pvag=0 delta=0.01 ngate=1e+030 dsub=0 cit=0.00114775 cdsc=0 
+ cdscd=1.99502e-005 cdscb=0 xpart=0 cgso=2.2653e-010 cgdo=2.2653e-010 cgbo=1e-013 cgsl=0 cgdl=0 ckappa=0.6 cf=0 clc=1e-007 cle=0.6 dlc=0 dwc=0 vfbcv=-0.826159 noff=1 voffcv=0 acde=0.5 moin=15 wln=1 wl=0 wwn=1 ww=0 wwl=0 lln=1 ll=0 lwn=1 lw=0 lwl=0 
+ llc=0 lwc=0 lwlc=0 wlc=0 wwc=0 wwlc=0 alpha0=0 alpha1=0 beta0=30 af=1.1021 kf=1.74179e-023 rsh=3 js=0.0001 jsw=0 cj=0.00150656 mj=0.403022 pb=0.790743 cjsw=1.18641e-010 mjsw=2 tref=27 prt=-149.998 ute=-0.950103 kt1=-0.257006 kt1l=0 kt2=-0.0222175 
+ ua1=1.29549e-010 ub1=-1.58953e-018 uc1=-4.01361e-011 at=-50000 xti=3 tcj=0.00075544 tcjsw=0.0017757 tpb=0.0016635 tpbsw=-0.0013729 elm=5 xl=0 xw=0 ldif=1e-007 hdif=2.7e-007 lmlt=1 wmlt=1 rd=0 rdc=0 rs=0 rsc=0 php=0.8 cjgate=2e-014 n=1 

.model rpl_rt r res=1 

.model mim_main c cap=1 tc1=2.5e-005 

.model vpnp1 pnp bf=1.3446 br=0.0179 is=3.75e-018 nf=1.069 nr=1.0037 isc=2.56e-017 ise=3.75e-018 nc=1.5 ne=2.083 vaf=485.868 var=10 ikf=0.000719 ikr=1.5 irb=9.9424 rb=85.468 re=0.1265 rc=1.686 cjc=9.99e-015 cje=1.089e-015 cjs=0 fc=0.75 mjc=0.39692 
+ mje=0.4409 mjs=0.5 vjc=0.677145 vje=0.9087 vjs=0.75 xcjc=0.5 cbcp=0 cbep=0 ccsp=0 itf=0.1 ptf=0 tf=1e-010 tr=0 vtf=10 xtf=1 af=1 kf=0 eg=1.224 xti=0.1825 tref=27 

.end
