module NOR2H(Q, X1, X2);
output Q;
input X1,X2;
nor(Q, X1,X2);
endmodule
