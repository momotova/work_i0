module NAND2H (Q, X1,X2);
    output Q;
    input X1,X2;
nand(Q, X1,X2);
endmodule
